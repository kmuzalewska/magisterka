library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => ("00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
1 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01"),
2 => ("01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
3 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
4 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00"),
5 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
6 => ("00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
7 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
8 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
9 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01")),
(
0 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00"),
1 => ("00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
2 => ("01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
3 => ("01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01"),
4 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01"),
5 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
6 => ("00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
7 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01"),
8 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00"),
9 => ("01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00")),
(
0 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11"),
1 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11"),
2 => ("01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00"),
3 => ("00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01"),
4 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
5 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11"),
6 => ("01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01"),
7 => ("00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
8 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00"),
9 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01")),
(
0 => ("01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01"),
1 => ("01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "11", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01"),
2 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "01", "11", "01", "01", "00"),
3 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
4 => ("00", "01", "00", "01", "01", "00", "11", "01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00"),
5 => ("00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "11", "00"),
6 => ("00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01"),
7 => ("00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00"),
8 => ("01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01"),
9 => ("01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00")),
(
0 => ("01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00"),
1 => ("00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "11", "11", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01"),
2 => ("01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "11", "00", "11"),
3 => ("00", "01", "00", "00", "11", "11", "00", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00"),
4 => ("01", "00", "00", "11", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01"),
5 => ("01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "11", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00"),
6 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "01", "01", "01", "11", "01", "11"),
7 => ("00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "11", "01", "11", "01", "00", "00", "01", "01", "01", "01"),
8 => ("01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "01", "01", "00"),
9 => ("01", "00", "01", "00", "00", "11", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "11", "01", "01", "01", "01", "01")),
(
0 => ("01", "00", "01", "01", "11", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "01", "11", "01", "01", "00", "01", "01"),
1 => ("01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "11", "11", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01"),
2 => ("00", "01", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11"),
3 => ("00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "11", "01", "00", "01", "01", "11", "01", "01", "11", "01"),
4 => ("01", "00", "00", "01", "00", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "11", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01"),
5 => ("01", "00", "01", "00", "11", "11", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00"),
6 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "11", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "00", "00", "00", "01", "00", "00"),
7 => ("01", "01", "00", "00", "11", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "11", "01", "11", "00"),
8 => ("00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "11", "00", "01", "01", "01", "01"),
9 => ("00", "11", "00", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00")),
(
0 => ("00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "11", "00", "00", "00", "00"),
1 => ("01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "11", "11", "01", "00", "11", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
2 => ("00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "00", "11", "01", "00", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "11", "11", "01", "00"),
3 => ("01", "01", "11", "00", "00", "01", "00", "00", "00", "11", "00", "11", "00", "11", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00"),
4 => ("01", "11", "00", "01", "11", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "11", "00", "01", "01", "11", "01"),
5 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "11", "00", "11", "01"),
6 => ("00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "00", "00", "11", "00", "11", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "01", "00", "11"),
7 => ("00", "11", "11", "01", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "11", "01", "00", "01", "00", "01"),
8 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "11", "11", "00", "00", "01", "00", "11", "11", "01", "00", "00", "00"),
9 => ("01", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "01", "00")),
(
0 => ("00", "11", "11", "11", "11", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "11"),
1 => ("01", "00", "11", "00", "11", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "11", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01"),
2 => ("01", "00", "00", "11", "00", "00", "01", "01", "01", "11", "00", "00", "11", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "00", "00", "11", "01", "00", "00", "01", "01"),
3 => ("00", "01", "01", "01", "00", "01", "01", "11", "01", "11", "01", "11", "00", "01", "00", "01", "01", "11", "11", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01"),
4 => ("01", "11", "00", "11", "11", "01", "00", "00", "00", "11", "00", "00", "01", "11", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01"),
5 => ("00", "00", "11", "00", "00", "01", "01", "11", "11", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
6 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "11", "11", "00", "11", "11", "11", "11", "00"),
7 => ("00", "11", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "11", "00", "11"),
8 => ("00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "11", "01", "01", "11", "11", "11", "11", "01", "00", "01", "01", "00"),
9 => ("01", "11", "00", "11", "00", "11", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "11", "00")),
(
0 => ("01", "01", "01", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00", "01", "01", "01", "01", "11", "01", "00"),
1 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "01", "00", "11", "01", "11", "01", "00", "01", "00", "11", "00", "01", "11", "11"),
2 => ("01", "01", "11", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "11", "00", "00", "01", "11", "11", "00", "00", "01", "01", "01", "01"),
3 => ("00", "01", "01", "00", "00", "00", "01", "11", "11", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "11", "11", "00", "01", "00", "00", "11", "00"),
4 => ("00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "11", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11"),
5 => ("01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "00", "00", "11", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "11", "00", "11", "00"),
6 => ("00", "11", "00", "11", "01", "00", "00", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "00", "01", "00", "11", "01"),
7 => ("00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "11", "01", "11", "11", "01", "01", "00", "01", "00", "11", "11", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
8 => ("01", "01", "00", "00", "11", "11", "11", "00", "01", "00", "01", "11", "11", "01", "01", "00", "01", "11", "11", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01"),
9 => ("01", "01", "11", "00", "01", "11", "11", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "11", "11", "01", "00", "01", "11", "01", "11", "00")),
(
0 => ("00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "11", "00", "11", "01", "00", "11", "01", "00", "11", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11"),
1 => ("00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "11", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "11", "00"),
2 => ("01", "01", "01", "11", "11", "11", "00", "01", "00", "01", "01", "00", "11", "00", "11", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "11", "01", "00", "00"),
3 => ("01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "11", "01", "01", "11", "01", "11", "01", "00", "11", "01", "11", "00", "00"),
4 => ("00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "11", "11", "00", "00", "01", "00", "11", "01", "01", "11", "00", "01", "11", "01", "00", "01", "01", "00", "11", "01", "00", "11"),
5 => ("00", "00", "01", "00", "00", "11", "00", "01", "11", "00", "11", "00", "00", "11", "01", "11", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "11", "11", "00"),
6 => ("01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "11", "11", "11", "01", "11", "00", "01", "00", "11", "01", "00", "11", "01", "01", "00", "01", "11", "00", "00", "00", "00"),
7 => ("00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "11", "11", "11", "11", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "11", "11"),
8 => ("01", "11", "00", "00", "00", "00", "11", "00", "11", "00", "01", "01", "00", "00", "11", "11", "01", "00", "00", "11", "01", "01", "11", "00", "01", "00", "01", "11", "01", "11", "01", "00"),
9 => ("00", "00", "00", "01", "01", "01", "11", "01", "11", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00", "11", "11", "11", "11", "01", "00", "01")));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;