library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => ("01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
1 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01"),
2 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
3 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
4 => ("01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
5 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
6 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
7 => ("00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00"),
8 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
9 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
others => (others =>"00")),
(
0 => ("00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01"),
1 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
2 => ("00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
3 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
4 => ("00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "00"),
5 => ("00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00"),
6 => ("00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
7 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01"),
8 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00"),
9 => ("01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
10 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
11 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00"),
12 => ("01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
13 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
14 => ("01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
15 => ("00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00"),
16 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01"),
17 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
18 => ("01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
19 => ("00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00"),
20 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00"),
21 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
22 => ("00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
23 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00"),
24 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
25 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00"),
26 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
27 => ("00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
28 => ("00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01"),
29 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
30 => ("01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01"),
31 => ("00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
32 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01"),
33 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00"),
34 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00"),
35 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
36 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00"),
37 => ("01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01"),
38 => ("00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
39 => ("01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
40 => ("01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
41 => ("01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00"),
42 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
43 => ("00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00"),
44 => ("00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01"),
45 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
46 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
47 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01"),
48 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00"),
49 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01"),
50 => ("00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
51 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01"),
52 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
53 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00"),
54 => ("01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01"),
55 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01"),
56 => ("00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01"),
57 => ("00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01"),
58 => ("00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
59 => ("00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01"),
60 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
61 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
62 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
63 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11"),
64 => ("01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00"),
65 => ("01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
66 => ("00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
67 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00"),
68 => ("01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01"),
69 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01"),
70 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00"),
71 => ("01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
72 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00"),
73 => ("00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
74 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00"),
75 => ("01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01"),
76 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
77 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
78 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
79 => ("00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
80 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00"),
81 => ("00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
82 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00"),
83 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
84 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00"),
85 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
86 => ("00", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
87 => ("01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
88 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
89 => ("00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
90 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00"),
91 => ("00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00"),
92 => ("00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00"),
93 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01"),
94 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00"),
95 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00"),
96 => ("00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
97 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01"),
98 => ("01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
99 => ("00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00"),
100 => ("01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
101 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00"),
102 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01"),
103 => ("00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
104 => ("01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00"),
105 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
106 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01"),
107 => ("01", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00"),
108 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
109 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
110 => ("00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00"),
111 => ("00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
112 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
113 => ("00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01"),
114 => ("01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
115 => ("00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
116 => ("01", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00"),
117 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
118 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
119 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
120 => ("01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00"),
121 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01"),
122 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01"),
123 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00"),
124 => ("01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01"),
125 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00"),
126 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01"),
127 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01"),
128 => ("00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
129 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00"),
130 => ("01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
131 => ("01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00"),
132 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00"),
133 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00"),
134 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01"),
135 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
136 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00"),
137 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
138 => ("01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
139 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
140 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
141 => ("01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
142 => ("00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
143 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
144 => ("01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
145 => ("01", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
146 => ("00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00"),
147 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11"),
148 => ("00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01"),
149 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01"),
150 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
151 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01"),
152 => ("01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01"),
153 => ("01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00"),
154 => ("01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
155 => ("00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
156 => ("00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
157 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01"),
158 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
159 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
160 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01"),
161 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00"),
162 => ("00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01"),
163 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01"),
164 => ("01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
165 => ("01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01"),
166 => ("00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00"),
167 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00"),
168 => ("01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01"),
169 => ("00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00"),
170 => ("00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
171 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01"),
172 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01"),
173 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
174 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11"),
175 => ("01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00"),
176 => ("01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01"),
177 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00"),
178 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01"),
179 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
180 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11"),
181 => ("00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
182 => ("00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00"),
183 => ("00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01"),
184 => ("01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
185 => ("00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00"),
186 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01"),
187 => ("01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00"),
188 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
189 => ("00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
190 => ("01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01"),
191 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
192 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01"),
193 => ("00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
194 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00"),
195 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01"),
196 => ("00", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
197 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01"),
198 => ("01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
199 => ("01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00"),
200 => ("01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01"),
201 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
202 => ("01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
203 => ("01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00"),
204 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11"),
205 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01"),
206 => ("00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
207 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
208 => ("00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
209 => ("01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
210 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "11"),
211 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00"),
212 => ("00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01"),
213 => ("01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
214 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
215 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01"),
216 => ("01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "01"),
217 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
218 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
219 => ("01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00"),
220 => ("00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01"),
221 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01"),
222 => ("01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00"),
223 => ("01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01"),
224 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01"),
225 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01"),
226 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01"),
227 => ("00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
228 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
229 => ("00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01"),
230 => ("01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01"),
231 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01"),
232 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00"),
233 => ("01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01"),
234 => ("00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01"),
235 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01"),
236 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
237 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
238 => ("01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00"),
239 => ("01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
240 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11"),
241 => ("00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
242 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
243 => ("01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
244 => ("01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00"),
245 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
246 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01"),
247 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00"),
248 => ("01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
249 => ("00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
250 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
251 => ("00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01"),
252 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01"),
253 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
254 => ("00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
255 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
256 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01"),
257 => ("01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
258 => ("00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
259 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00"),
260 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01"),
261 => ("01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
262 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
263 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
264 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01"),
265 => ("00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01"),
266 => ("01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01"),
267 => ("00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01"),
268 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01"),
269 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
270 => ("01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
271 => ("00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
272 => ("01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00"),
273 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01"),
274 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
275 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01"),
276 => ("01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00"),
277 => ("00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
278 => ("01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00"),
279 => ("01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
280 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
281 => ("00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
282 => ("00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
283 => ("00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
284 => ("00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01"),
285 => ("00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
286 => ("00", "01", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
287 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00"),
288 => ("01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
289 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00"),
290 => ("01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
291 => ("01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00"),
292 => ("00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
293 => ("00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01"),
294 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00"),
295 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
296 => ("00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
297 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00"),
298 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
299 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
300 => ("00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
301 => ("00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00"),
302 => ("00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01"),
303 => ("00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
304 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01"),
305 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00"),
306 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01"),
307 => ("01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00"),
308 => ("00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00"),
309 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
310 => ("00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00"),
311 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
312 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01"),
313 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
314 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11"),
315 => ("01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00"),
316 => ("00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
317 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01"),
318 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01"),
319 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01"),
320 => ("01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
321 => ("00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
322 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
323 => ("00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
324 => ("01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
325 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
326 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01"),
327 => ("00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
328 => ("00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
329 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01"),
330 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01"),
331 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01"),
332 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01"),
333 => ("00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
334 => ("00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
335 => ("00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
336 => ("00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00"),
337 => ("01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
338 => ("01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01"),
339 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "00"),
340 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
341 => ("00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01"),
342 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
343 => ("00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11"),
344 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00"),
345 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
346 => ("00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11"),
347 => ("01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
348 => ("00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
349 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00"),
350 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00"),
351 => ("00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
352 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
353 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01"),
354 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00"),
355 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
356 => ("01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
357 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01"),
358 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01"),
359 => ("01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00"),
360 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00"),
361 => ("00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
362 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01"),
363 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01"),
364 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
365 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
366 => ("00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00"),
367 => ("00", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
368 => ("01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00"),
369 => ("01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01"),
370 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
371 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00"),
372 => ("00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
373 => ("00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01"),
374 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11"),
375 => ("00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
376 => ("01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01"),
377 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
378 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01"),
379 => ("01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
380 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
381 => ("00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01"),
382 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01"),
383 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
384 => ("00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
385 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
386 => ("01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
387 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
388 => ("01", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
389 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
390 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00"),
391 => ("01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
392 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00"),
393 => ("00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00"),
394 => ("01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
395 => ("01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00"),
396 => ("00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00"),
397 => ("00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
398 => ("00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11"),
399 => ("01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
400 => ("00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01"),
401 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01"),
402 => ("00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00"),
403 => ("00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
404 => ("01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01"),
405 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01"),
406 => ("00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
407 => ("01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
408 => ("00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
409 => ("00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01"),
410 => ("00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
411 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11"),
412 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00"),
413 => ("01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01"),
414 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00"),
415 => ("00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00"),
416 => ("01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00"),
417 => ("01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
418 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
419 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
420 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00"),
421 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00"),
422 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00"),
423 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01"),
424 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01"),
425 => ("01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01"),
426 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
427 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
428 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
429 => ("01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01"),
430 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
431 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11"),
432 => ("01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
433 => ("01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
434 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
435 => ("01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
436 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
437 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
438 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00"),
439 => ("00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
440 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
441 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00"),
442 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00"),
443 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01"),
444 => ("01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01"),
445 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00"),
446 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
447 => ("00", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01"),
448 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00"),
449 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01"),
450 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00"),
451 => ("00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00"),
452 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01"),
453 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
454 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
455 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
456 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00"),
457 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
458 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
459 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01"),
460 => ("01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
461 => ("01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00"),
462 => ("01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
463 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "00"),
464 => ("01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
465 => ("01", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
466 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00"),
467 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
468 => ("01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
469 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00"),
470 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
471 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
472 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01"),
473 => ("01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01"),
474 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01"),
475 => ("01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
476 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01"),
477 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01"),
478 => ("01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00"),
479 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "01"),
480 => ("00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01"),
481 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00"),
482 => ("01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
483 => ("00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
484 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00"),
485 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
486 => ("01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01"),
487 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01"),
488 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01"),
489 => ("01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
490 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01"),
491 => ("01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
492 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
493 => ("01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01"),
494 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00"),
495 => ("01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
496 => ("01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00"),
497 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
498 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
499 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
500 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00"),
501 => ("00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01"),
502 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "01"),
503 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00"),
504 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01"),
505 => ("00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01"),
506 => ("00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00"),
507 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01"),
508 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11"),
509 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
510 => ("00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
511 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01"),
512 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
513 => ("01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
514 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
515 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
516 => ("01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00"),
517 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
518 => ("00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00"),
519 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11"),
520 => ("00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01"),
521 => ("01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00"),
522 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
523 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01"),
524 => ("00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11"),
525 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00"),
526 => ("01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
527 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
528 => ("00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01"),
529 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
530 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "00"),
531 => ("00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01"),
532 => ("01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01"),
533 => ("01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01"),
534 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
535 => ("01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
536 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01"),
537 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00"),
538 => ("01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01"),
539 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00"),
540 => ("00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
541 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01"),
542 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01"),
543 => ("01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
544 => ("00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01"),
545 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
546 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01"),
547 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01"),
548 => ("00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
549 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01"),
550 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "00"),
551 => ("01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00"),
552 => ("01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
553 => ("00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01"),
554 => ("01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
555 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00"),
556 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00"),
557 => ("01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
558 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
559 => ("01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
560 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "01", "00", "01"),
561 => ("00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
562 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01"),
563 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
564 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
565 => ("01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
566 => ("01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00"),
567 => ("01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
568 => ("00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
569 => ("00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
570 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00"),
571 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01"),
572 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
573 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01"),
574 => ("00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
575 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00"),
576 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
577 => ("01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
578 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
579 => ("01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01"),
580 => ("00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01"),
581 => ("00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
582 => ("01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01"),
583 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
584 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
585 => ("01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01"),
586 => ("01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
587 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
588 => ("01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01"),
589 => ("00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
590 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
591 => ("01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00"),
592 => ("01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
593 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "00"),
594 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01"),
595 => ("00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01"),
596 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "00"),
597 => ("01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00"),
598 => ("00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
599 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01"),
600 => ("00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00"),
601 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01"),
602 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00"),
603 => ("00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
604 => ("01", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
605 => ("00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
606 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "00"),
607 => ("01", "00", "01", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
608 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
609 => ("00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
610 => ("00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
611 => ("00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00"),
612 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
613 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01"),
614 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01"),
615 => ("01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01"),
616 => ("00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01"),
617 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00"),
618 => ("00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00"),
619 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01"),
620 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00"),
621 => ("00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01"),
622 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01"),
623 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
624 => ("01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
625 => ("01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00"),
626 => ("00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
627 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
628 => ("01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
629 => ("01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
630 => ("00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
631 => ("01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00"),
632 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00"),
633 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01"),
634 => ("00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
635 => ("00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
636 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00"),
637 => ("00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
638 => ("00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
639 => ("00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01"),
640 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01"),
641 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01"),
642 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00"),
643 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
644 => ("00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
645 => ("01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00"),
646 => ("00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
647 => ("00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01"),
648 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
649 => ("00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00"),
650 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01"),
651 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
652 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00"),
653 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
654 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01"),
655 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
656 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00"),
657 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
658 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
659 => ("00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00"),
660 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00"),
661 => ("00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
662 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
663 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
664 => ("00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00"),
665 => ("01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
666 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
667 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
668 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
669 => ("00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01"),
670 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01"),
671 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11"),
672 => ("00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
673 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
674 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00"),
675 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
676 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00"),
677 => ("01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
678 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00"),
679 => ("00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01"),
680 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
681 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01"),
682 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
683 => ("00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01"),
684 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
685 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
686 => ("00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01"),
687 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
688 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01"),
689 => ("01", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
690 => ("00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
691 => ("01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
692 => ("00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00"),
693 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11"),
694 => ("00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
695 => ("00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00"),
696 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
697 => ("01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01"),
698 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00"),
699 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
700 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00"),
701 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00"),
702 => ("01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00"),
703 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
704 => ("01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11"),
705 => ("01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00"),
706 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01"),
707 => ("00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
708 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
709 => ("00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01"),
710 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
711 => ("00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
712 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01"),
713 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
714 => ("01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01"),
715 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
716 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
717 => ("01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00"),
718 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01"),
719 => ("01", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00"),
720 => ("01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
721 => ("00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
722 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
723 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11"),
724 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
725 => ("01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
726 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01"),
727 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
728 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
729 => ("00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00"),
730 => ("01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01"),
731 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00"),
732 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
733 => ("00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01"),
734 => ("01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01"),
735 => ("01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01"),
736 => ("01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01"),
737 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00"),
738 => ("00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
739 => ("00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
740 => ("01", "00", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
741 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01"),
742 => ("01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
743 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01"),
744 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
745 => ("01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
746 => ("01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00"),
747 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01"),
748 => ("00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01"),
749 => ("01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
750 => ("01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01"),
751 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00"),
752 => ("00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00"),
753 => ("01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
754 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
755 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01"),
756 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01"),
757 => ("00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01"),
758 => ("00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
759 => ("01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
760 => ("01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01"),
761 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
762 => ("00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00"),
763 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01"),
764 => ("01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
765 => ("01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
766 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01"),
767 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00"),
768 => ("01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00"),
769 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01"),
770 => ("00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
771 => ("00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01"),
772 => ("00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00"),
773 => ("00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
774 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00"),
775 => ("01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00"),
776 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00"),
777 => ("01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
778 => ("00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
779 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
780 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00"),
781 => ("00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00"),
782 => ("01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
783 => ("00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01"),
784 => ("01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00"),
785 => ("01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01"),
786 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00"),
787 => ("00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
788 => ("00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00"),
789 => ("00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
790 => ("00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
791 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00"),
792 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
793 => ("01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
794 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "11"),
795 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11"),
796 => ("00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01"),
797 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01"),
798 => ("01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
799 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
800 => ("01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
801 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
802 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01"),
803 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00"),
804 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
805 => ("00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
806 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00"),
807 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01"),
808 => ("00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00"),
809 => ("01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00"),
810 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
811 => ("01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01"),
812 => ("01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
813 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00"),
814 => ("01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01"),
815 => ("00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00"),
816 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
817 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01"),
818 => ("01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00"),
819 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01"),
820 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
821 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00"),
822 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
823 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
824 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01"),
825 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00"),
826 => ("00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
827 => ("01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
828 => ("00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00"),
829 => ("00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
830 => ("00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
831 => ("01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
832 => ("01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
833 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00"),
834 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01"),
835 => ("01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01"),
836 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
837 => ("00", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
838 => ("01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
839 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
840 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
841 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01"),
842 => ("01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01"),
843 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00"),
844 => ("01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00"),
845 => ("00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
846 => ("00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
847 => ("00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
848 => ("00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
849 => ("01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01"),
850 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
851 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
852 => ("00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
853 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
854 => ("01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00"),
855 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00"),
856 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01"),
857 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01"),
858 => ("01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01"),
859 => ("00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
860 => ("00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00"),
861 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
862 => ("01", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
863 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
864 => ("01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
865 => ("00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
866 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01"),
867 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
868 => ("00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
869 => ("01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
870 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
871 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
872 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
873 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
874 => ("01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00"),
875 => ("01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01"),
876 => ("01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00"),
877 => ("00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
878 => ("00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00"),
879 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
880 => ("01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
881 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01"),
882 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
883 => ("01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01"),
884 => ("01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
885 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
886 => ("00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00"),
887 => ("00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
888 => ("01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01"),
889 => ("00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01"),
890 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01"),
891 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
892 => ("01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01"),
893 => ("01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00"),
894 => ("01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00"),
895 => ("01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01"),
896 => ("00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01"),
897 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
898 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
899 => ("00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00"),
900 => ("00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01"),
901 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01"),
902 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01"),
903 => ("00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00"),
904 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
905 => ("00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
906 => ("00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01"),
907 => ("00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01"),
908 => ("01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00"),
909 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
910 => ("00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
911 => ("00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
912 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00"),
913 => ("01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
914 => ("01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"),
915 => ("01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
916 => ("00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01"),
917 => ("01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
918 => ("01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
919 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
920 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01"),
921 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "00"),
922 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00"),
923 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
924 => ("01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
925 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00"),
926 => ("01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00"),
927 => ("01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
928 => ("00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11"),
929 => ("00", "01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
930 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
931 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00"),
932 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
933 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00"),
934 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00"),
935 => ("01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00"),
936 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01"),
937 => ("00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
938 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
939 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01"),
940 => ("01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
941 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
942 => ("01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01"),
943 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
944 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00"),
945 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
946 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00"),
947 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
948 => ("00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
949 => ("01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
950 => ("00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00"),
951 => ("00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00"),
952 => ("00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00"),
953 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00"),
954 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00"),
955 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01"),
956 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
957 => ("01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00"),
958 => ("00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00"),
959 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00"),
960 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01"),
961 => ("01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00"),
962 => ("00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
963 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00"),
964 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00"),
965 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
966 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00"),
967 => ("00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
968 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00"),
969 => ("01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00"),
970 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
971 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01"),
972 => ("01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00"),
973 => ("00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00"),
974 => ("01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00"),
975 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01"),
976 => ("01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01"),
977 => ("00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00"),
978 => ("01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
979 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
980 => ("01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
981 => ("00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
982 => ("01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
983 => ("01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
984 => ("00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
985 => ("00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00"),
986 => ("01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
987 => ("00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01"),
988 => ("00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00"),
989 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00"),
990 => ("01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
991 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01"),
992 => ("01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01"),
993 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
994 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00"),
995 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
996 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01"),
997 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00"),
998 => ("01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00"),
999 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01")),
(
0 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01"),
1 => ("00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11"),
2 => ("01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01"),
3 => ("00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01"),
4 => ("01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00"),
5 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
6 => ("00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00"),
7 => ("00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00"),
8 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01"),
9 => ("01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01"),
others => (others =>"00")),
(
0 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "11", "01", "11", "00", "00"),
1 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "01", "11", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "00"),
2 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00"),
3 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01"),
4 => ("01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01"),
5 => ("00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
6 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01"),
7 => ("01", "01", "01", "00", "11", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
8 => ("01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00"),
9 => ("00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
others => (others =>"00")),
(
0 => ("00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "11", "01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
1 => ("00", "11", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00"),
2 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "11", "00", "00", "01", "00", "01", "11"),
3 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "11", "00", "00", "00", "01", "01", "11", "01"),
4 => ("00", "11", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "11", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01"),
5 => ("01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "11", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00"),
6 => ("01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "11"),
7 => ("00", "01", "00", "11", "01", "00", "11", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01"),
8 => ("01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "11", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00"),
9 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00"),
others => (others =>"00")),
(
0 => ("01", "00", "00", "01", "00", "11", "01", "00", "11", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "11", "00", "00"),
1 => ("00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "00", "01", "11", "00", "01", "00", "01", "01", "11", "11", "01", "00", "01", "00", "01"),
2 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "11", "00", "01", "11", "00", "11"),
3 => ("01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "11", "01", "11"),
4 => ("00", "00", "11", "01", "01", "01", "11", "11", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
5 => ("00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "11", "00", "00", "01", "11"),
6 => ("00", "11", "00", "11", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
7 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01"),
8 => ("01", "00", "01", "00", "00", "00", "01", "11", "00", "11", "01", "01", "01", "11", "00", "11", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
9 => ("00", "11", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "11", "01", "00", "01", "01", "01"),
others => (others =>"00")),
(
0 => ("01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "11", "11", "00", "00", "01", "11"),
1 => ("00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "11", "01", "01", "00", "11", "11", "01", "00", "00", "11", "00", "11", "01", "01", "01", "01", "01", "01"),
2 => ("00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "11", "00", "11", "01", "01"),
3 => ("01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "11", "11", "00", "00", "01", "11", "01", "01", "01", "00"),
4 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "11", "11", "11", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11"),
5 => ("01", "00", "11", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "01", "01", "01", "01"),
6 => ("00", "11", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01"),
7 => ("00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "11", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "11"),
8 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "11", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "11", "11", "11", "01", "00", "00", "01"),
9 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "11", "11", "11", "11", "00", "01"),
others => (others =>"00")),
(
0 => ("00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "01", "11", "11", "01", "00", "01", "01", "11", "11", "01", "00", "00", "01"),
1 => ("00", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "11", "01", "11", "01", "00", "11", "00", "01", "11", "00", "00", "01", "01"),
2 => ("01", "01", "11", "11", "01", "11", "11", "11", "00", "00", "11", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
3 => ("01", "01", "01", "00", "11", "11", "00", "01", "01", "00", "01", "01", "00", "11", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "11"),
4 => ("00", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00", "11", "00", "00", "11", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "11", "11", "01", "00", "00"),
5 => ("00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "11", "01", "00", "11", "11", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01"),
6 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "11", "00", "01", "00", "00", "11", "01", "00", "11", "00", "11", "00", "00", "01", "00", "01", "00", "01", "11", "00", "11"),
7 => ("01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "11", "01", "01", "00", "11", "00", "01", "01", "11", "01", "01", "00", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00"),
8 => ("01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "11", "11", "01", "00", "00", "11", "00", "01", "11", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11"),
9 => ("01", "11", "00", "00", "11", "01", "11", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "11", "01", "01", "01"),
others => (others =>"00")),
(
0 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "11", "11", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01", "11"),
1 => ("00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "11", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01"),
2 => ("00", "00", "11", "00", "11", "00", "11", "00", "01", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "11", "00", "01", "00"),
3 => ("01", "00", "00", "11", "00", "01", "11", "11", "01", "00", "00", "01", "01", "01", "01", "00", "11", "11", "00", "01", "00", "01", "01", "11", "00", "11", "01", "01", "00", "00", "00", "00"),
4 => ("00", "00", "00", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "00", "11", "01", "11", "00", "01", "01", "11", "01", "01", "01", "01", "11", "01", "01", "01", "11", "01"),
5 => ("01", "00", "00", "00", "00", "11", "01", "11", "11", "01", "01", "00", "00", "01", "00", "01", "00", "11", "11", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01"),
6 => ("01", "00", "00", "01", "11", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "11", "01", "00", "00", "11", "00", "00", "01", "00", "01", "11", "01", "00", "00", "11", "00", "00"),
7 => ("01", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01", "11", "00", "11", "11", "00", "01", "11", "00", "11", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01"),
8 => ("00", "11", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "11", "00", "00", "00", "11", "11", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "11", "00", "01", "01"),
9 => ("01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "11", "01", "11", "00", "00", "11", "00", "00", "01", "11", "00", "01", "01", "01"),
others => (others =>"00")),
(
0 => ("00", "00", "00", "11", "00", "11", "01", "11", "00", "01", "01", "00", "00", "11", "00", "01", "01", "11", "00", "11", "01", "11", "00", "00", "01", "01", "01", "11", "01", "01", "11", "01"),
1 => ("00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "11", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "00", "00", "11", "11", "01", "01", "11", "11", "11"),
2 => ("00", "00", "11", "11", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "11", "00", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
3 => ("01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "11", "00", "00", "01", "11", "11", "11", "01", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "01", "01", "11", "00"),
4 => ("00", "01", "00", "00", "01", "11", "00", "00", "11", "01", "11", "00", "00", "00", "11", "00", "11", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "00", "01", "00", "00", "11"),
5 => ("00", "01", "01", "11", "11", "00", "01", "11", "01", "01", "11", "11", "11", "01", "00", "11", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01"),
6 => ("00", "01", "11", "01", "11", "00", "11", "11", "11", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01"),
7 => ("01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "11"),
8 => ("01", "11", "00", "11", "11", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "11", "11", "01", "01", "01", "11", "01", "00", "11", "00", "00", "00", "01", "00"),
9 => ("00", "00", "11", "01", "01", "00", "01", "11", "01", "00", "01", "00", "11", "11", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "11", "00", "11", "00", "00"),
others => (others =>"00")));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;