library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
1 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01"),
2 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00"),
3 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00"),
4 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00"),
5 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
6 => ("01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01"),
7 => ("01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
8 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
9 => ("01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00"),
others => (others =>"00")),
(
0 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00"),
1 => ("01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01"),
2 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00"),
3 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01"),
4 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
5 => ("01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01"),
6 => ("01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01"),
7 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
8 => ("01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
9 => ("01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01"),
10 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
11 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01"),
12 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
13 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00"),
14 => ("00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
15 => ("00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
16 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00"),
17 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
18 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
19 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01"),
20 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11"),
21 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01"),
22 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00"),
23 => ("00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01"),
24 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
25 => ("01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00"),
26 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01"),
27 => ("00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01"),
28 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
29 => ("00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
30 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01"),
31 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
32 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11"),
33 => ("00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
34 => ("00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01"),
35 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
36 => ("00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
37 => ("01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00"),
38 => ("01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01"),
39 => ("01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
40 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
41 => ("01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00"),
42 => ("00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
43 => ("00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
44 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "01", "00"),
45 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
46 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "00"),
47 => ("01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
48 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00"),
49 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00"),
50 => ("01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
51 => ("00", "00", "01", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
52 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01"),
53 => ("01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
54 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00"),
55 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01"),
56 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00"),
57 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01"),
58 => ("01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
59 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00"),
60 => ("00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01"),
61 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00"),
62 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00"),
63 => ("00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
64 => ("00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
65 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01"),
66 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01"),
67 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01"),
68 => ("01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01"),
69 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01"),
70 => ("01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01"),
71 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01"),
72 => ("01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01"),
73 => ("01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
74 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11"),
75 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01"),
76 => ("01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
77 => ("01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01"),
78 => ("01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
79 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
80 => ("01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01"),
81 => ("00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01"),
82 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
83 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
84 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
85 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
86 => ("01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01"),
87 => ("01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01"),
88 => ("01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
89 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01"),
90 => ("01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
91 => ("00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01"),
92 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
93 => ("00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
94 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00"),
95 => ("01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
96 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
97 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00"),
98 => ("00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00"),
99 => ("00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01"),
100 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00"),
101 => ("00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
102 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00"),
103 => ("01", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
104 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
105 => ("01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00"),
106 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00"),
107 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
108 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
109 => ("00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00"),
110 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01"),
111 => ("01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00"),
112 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00"),
113 => ("01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
114 => ("00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01"),
115 => ("01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00"),
116 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01"),
117 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
118 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01"),
119 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00"),
120 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01"),
121 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
122 => ("00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
123 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00"),
124 => ("00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
125 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00"),
126 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
127 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
128 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01"),
129 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
130 => ("01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00"),
131 => ("01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00"),
132 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01"),
133 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
134 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00"),
135 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
136 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
137 => ("00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
138 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
139 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00"),
140 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01"),
141 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01"),
142 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
143 => ("01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01"),
144 => ("01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
145 => ("01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
146 => ("01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
147 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01"),
148 => ("01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
149 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
150 => ("00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
151 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
152 => ("01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01"),
153 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00"),
154 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "01", "01"),
155 => ("00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00"),
156 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00"),
157 => ("00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
158 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01"),
159 => ("01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00"),
160 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
161 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00"),
162 => ("01", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01"),
163 => ("00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
164 => ("01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00"),
165 => ("01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00"),
166 => ("00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
167 => ("01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
168 => ("01", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
169 => ("01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
170 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00"),
171 => ("00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01"),
172 => ("00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00"),
173 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01"),
174 => ("01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00"),
175 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
176 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01"),
177 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00"),
178 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00"),
179 => ("01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00"),
180 => ("00", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
181 => ("00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00"),
182 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00"),
183 => ("00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01"),
184 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00"),
185 => ("00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
186 => ("00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
187 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
188 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
189 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01"),
190 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01"),
191 => ("00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
192 => ("01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00"),
193 => ("00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00"),
194 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
195 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
196 => ("01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00"),
197 => ("01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00"),
198 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01"),
199 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00"),
200 => ("01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01"),
201 => ("00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00"),
202 => ("00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00"),
203 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00"),
204 => ("00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
205 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00"),
206 => ("00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
207 => ("00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
208 => ("01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01"),
209 => ("01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01"),
210 => ("01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01"),
211 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01"),
212 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
213 => ("00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
214 => ("00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01"),
215 => ("01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "11", "01"),
216 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
217 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
218 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01"),
219 => ("00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
220 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00"),
221 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01"),
222 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
223 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00"),
224 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
225 => ("01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
226 => ("00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01"),
227 => ("01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
228 => ("00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01"),
229 => ("00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
230 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01"),
231 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
232 => ("01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
233 => ("01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01"),
234 => ("00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11"),
235 => ("01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
236 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
237 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00"),
238 => ("01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
239 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
240 => ("00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00"),
241 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
242 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00"),
243 => ("01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01"),
244 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01"),
245 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
246 => ("01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00"),
247 => ("00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
248 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01"),
249 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00"),
250 => ("00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00"),
251 => ("01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
252 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00"),
253 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
254 => ("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
255 => ("01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
256 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01"),
257 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00"),
258 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01"),
259 => ("01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
260 => ("00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
261 => ("01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01"),
262 => ("01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00"),
263 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
264 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01"),
265 => ("01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
266 => ("01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00"),
267 => ("01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
268 => ("00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
269 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
270 => ("00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
271 => ("01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00"),
272 => ("00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
273 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
274 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
275 => ("00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
276 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "00"),
277 => ("01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01"),
278 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
279 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
280 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01"),
281 => ("01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00"),
282 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "01"),
283 => ("01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
284 => ("00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
285 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01"),
286 => ("01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
287 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00"),
288 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
289 => ("01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
290 => ("01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
291 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00"),
292 => ("01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
293 => ("01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
294 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01"),
295 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00"),
296 => ("01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01"),
297 => ("00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01"),
298 => ("00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00"),
299 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
300 => ("01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
301 => ("00", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00"),
302 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01"),
303 => ("01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
304 => ("01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11"),
305 => ("01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
306 => ("01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00"),
307 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00"),
308 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01"),
309 => ("00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
310 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00"),
311 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00"),
312 => ("01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01"),
313 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01"),
314 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
315 => ("00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
316 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00"),
317 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01"),
318 => ("01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
319 => ("01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
320 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01"),
321 => ("00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00"),
322 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
323 => ("00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
324 => ("01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01"),
325 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
326 => ("01", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01"),
327 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01"),
328 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00"),
329 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
330 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
331 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00"),
332 => ("01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01"),
333 => ("01", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
334 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01"),
335 => ("00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00"),
336 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00"),
337 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
338 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01"),
339 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
340 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
341 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01"),
342 => ("01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
343 => ("00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
344 => ("00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
345 => ("01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
346 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "01"),
347 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01"),
348 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11"),
349 => ("01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
350 => ("01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01"),
351 => ("00", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
352 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
353 => ("01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01"),
354 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01"),
355 => ("00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
356 => ("01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
357 => ("00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01"),
358 => ("01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01"),
359 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
360 => ("00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
361 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01"),
362 => ("01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
363 => ("00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00"),
364 => ("01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
365 => ("01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
366 => ("01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00"),
367 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "00"),
368 => ("00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00"),
369 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11"),
370 => ("01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01"),
371 => ("00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "00"),
372 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
373 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01"),
374 => ("01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01"),
375 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
376 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
377 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01"),
378 => ("01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
379 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01"),
380 => ("01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
381 => ("00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01"),
382 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00"),
383 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00"),
384 => ("01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00"),
385 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00"),
386 => ("01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
387 => ("00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00"),
388 => ("00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01"),
389 => ("01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
390 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00"),
391 => ("00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01"),
392 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00"),
393 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11"),
394 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00"),
395 => ("01", "00", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
396 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
397 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "01"),
398 => ("00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00"),
399 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00")),
(
0 => ("01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00"),
1 => ("00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01"),
2 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
3 => ("01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00"),
4 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00"),
5 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11"),
6 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11"),
7 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11"),
8 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00"),
9 => ("01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01"),
others => (others =>"00")),
(
0 => ("00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00"),
1 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00"),
2 => ("00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11"),
3 => ("01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01"),
4 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "11", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01"),
5 => ("00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "01"),
6 => ("00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "11", "01", "00", "01", "00"),
7 => ("00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00"),
8 => ("00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01"),
9 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "11", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
others => (others =>"00")),
(
0 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "11"),
1 => ("00", "00", "01", "00", "01", "11", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "11"),
2 => ("00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "11", "00", "00", "01", "00", "00"),
3 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "11", "11", "01", "01"),
4 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "11", "01", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01"),
5 => ("01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "11", "11", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
6 => ("00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11"),
7 => ("00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "11"),
8 => ("01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "11", "01"),
9 => ("01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00"),
others => (others =>"00")),
(
0 => ("01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00"),
1 => ("00", "11", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01"),
2 => ("00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "00", "01", "11", "01", "00", "01"),
3 => ("00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "11", "00", "11", "01", "00"),
4 => ("01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "11", "00", "01", "00", "11", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00"),
5 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "11", "01", "01", "01", "00", "11", "01", "11", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00"),
6 => ("01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "11", "01"),
7 => ("01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "11", "00", "00", "11", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01"),
8 => ("01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "00", "11", "00", "11", "01", "01", "01"),
9 => ("01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "11"),
others => (others =>"00")),
(
0 => ("00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "00", "01", "11", "01", "01", "11", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00"),
1 => ("01", "01", "11", "01", "01", "01", "00", "11", "01", "01", "11", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "01", "01", "00", "01", "00", "01"),
2 => ("01", "11", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "11", "01", "00", "00"),
3 => ("00", "00", "00", "01", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "11", "00", "00", "11", "00", "01", "00"),
4 => ("00", "01", "11", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "11", "11", "00", "00", "01", "00", "00", "01", "11", "11", "01", "01", "00", "01", "01", "00"),
5 => ("01", "11", "01", "01", "00", "11", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01"),
6 => ("01", "01", "11", "01", "00", "01", "00", "01", "00", "11", "11", "00", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00"),
7 => ("01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "11", "00", "00", "00", "00", "11", "11", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "11"),
8 => ("01", "00", "11", "01", "01", "00", "11", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "11", "00", "00", "01", "01"),
9 => ("01", "00", "00", "00", "00", "01", "11", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "11", "00", "01", "01"),
others => (others =>"00")),
(
0 => ("00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "11", "00", "01", "11", "01", "01", "00", "11", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "11", "01"),
1 => ("00", "00", "01", "00", "00", "01", "00", "11", "11", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "11", "00", "00", "00", "00", "01", "00", "11", "11", "11", "01", "00", "01"),
2 => ("01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "11", "01", "00", "11", "00", "00", "11", "01", "00", "01"),
3 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "11", "11", "00", "01", "01", "11", "00", "01", "01", "11", "11", "11"),
4 => ("01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "01", "00", "01", "11", "11", "00", "11", "00", "01", "01", "11", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00"),
5 => ("01", "01", "00", "01", "00", "00", "11", "11", "11", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "01"),
6 => ("01", "00", "11", "01", "11", "00", "11", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01"),
7 => ("01", "11", "00", "01", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "11", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00"),
8 => ("01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "00", "11", "11", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "11"),
9 => ("00", "01", "01", "11", "11", "11", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
others => (others =>"00")),
(
0 => ("01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "11", "11", "01", "00", "01", "11", "01", "11", "01", "00", "01", "11", "00", "11", "01", "01", "01", "00", "01"),
1 => ("00", "11", "00", "11", "00", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11"),
2 => ("00", "11", "01", "01", "00", "11", "01", "11", "01", "01", "00", "00", "11", "00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "00", "11", "11", "01"),
3 => ("01", "01", "11", "11", "01", "01", "00", "00", "01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01"),
4 => ("01", "01", "00", "00", "11", "01", "11", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "11", "11", "00", "01", "11", "11", "00", "00", "01", "00", "01", "00", "11", "01", "00"),
5 => ("01", "11", "01", "11", "01", "11", "00", "00", "00", "01", "11", "01", "11", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "11", "01"),
6 => ("00", "11", "00", "01", "00", "00", "11", "11", "01", "11", "11", "00", "01", "11", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
7 => ("01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "11", "00", "11", "01", "00", "00", "01", "00", "11", "00", "00", "11", "11", "01", "00", "11", "01", "00", "00"),
8 => ("01", "11", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "01", "11", "11"),
9 => ("00", "11", "01", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "11", "11", "11", "00", "00", "01", "01", "00", "00", "00", "00", "11"),
others => (others =>"00")),
(
0 => ("01", "11", "01", "11", "11", "00", "00", "00", "00", "01", "00", "01", "11", "00", "11", "01", "01", "01", "11", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11"),
1 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "11", "11", "01", "11", "00", "01", "11", "01", "00", "00", "11", "11", "01", "01", "01"),
2 => ("01", "11", "11", "00", "01", "01", "11", "01", "11", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "11", "11", "01", "11", "11", "01", "00", "01", "01", "01", "00", "01"),
3 => ("01", "01", "00", "00", "11", "01", "00", "11", "00", "01", "01", "11", "00", "00", "00", "01", "11", "00", "00", "00", "01", "11", "01", "00", "11", "11", "00", "11", "01", "01", "11", "00"),
4 => ("01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "11", "11", "01", "11", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00", "01", "11", "11", "01"),
5 => ("00", "00", "01", "11", "11", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "11", "11", "01", "11", "00"),
6 => ("01", "01", "11", "00", "00", "11", "11", "01", "00", "00", "00", "00", "11", "00", "01", "00", "01", "11", "01", "11", "01", "00", "11", "01", "01", "00", "11", "00", "01", "11", "01", "00"),
7 => ("01", "01", "00", "01", "00", "11", "11", "01", "01", "11", "00", "11", "00", "00", "11", "11", "11", "11", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
8 => ("00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00", "11", "11", "01", "00", "01"),
9 => ("01", "11", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "01", "00", "00", "01", "00", "11", "01", "11", "11", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "11"),
others => (others =>"00")));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;