library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => "01011011000101010101011001110010",
1 => "01101110111001010101100101110000",
2 => "10110100100011011010100111100110",
3 => "10000111100010111010001111000010",
4 => "11000101100011110010000110101000",
5 => "10110100001111010110001011011100",
6 => "01010100010000100000000101100000",
7 => "11100001010101100101110110000011",
8 => "00111100101000101110111110100001",
9 => "11011000101011100110000101011100",
10 => "10000000001110100010101001010001",
11 => "01010010000100010000101001110010",
12 => "10101111110101000000101011000101",
13 => "10001100110101101010011000000110",
14 => "00011010000111111100010010000001",
15 => "00010111001010010001110010101011",
16 => "10011110110010011000110000001110",
17 => "11011001100000011001001001111000",
18 => "01110011111010000100100101010101",
19 => "10100001010100011110111100010001",
20 => "10110000000000011011111100011110",
21 => "00111101000010010111111011100110",
22 => "10000100110110110110101011000100",
23 => "11011010001101110001110111110110",
24 => "10000110100010000001110011110000",
25 => "11010010011000000100011101010011",
26 => "01111001110011011011110110000001",
27 => "10100110111111110101111001010101",
28 => "10100111000100001100000110110010",
29 => "11001010001011000101010000001110",
30 => "11111001000010111001011001011110",
31 => "01011001110111100111101101001110",
32 => "10101011001110100100111101101100",
33 => "01011110001011101101000110110001",
34 => "00101111100101100101110100111111",
35 => "00010111010111110111101101100111",
36 => "10111001101100000001101010001110",
37 => "10001110001100010110100000111001",
38 => "00100011101101001010011011000111",
39 => "11111010110000000001111101011011",
40 => "10101000010010001110011010000011",
41 => "01110110100111010100001100011101",
42 => "00110011010101110110000001011101",
43 => "11011111010111000001100100101101",
44 => "00111000001101001111011110001110",
45 => "11110101100001000101101111010000",
46 => "00111010011011000000001111010110",
47 => "01010100111110100011100000100110",
48 => "11100000011001111000011000111111",
49 => "00110001100000000001000000011111",
50 => "00011101011001101110110000111101",
51 => "00110101010110011010011000100100",
52 => "01101010011101111011011001100100",
53 => "01101110001001111011011001011101",
54 => "00100000010101001000111111101011",
55 => "01101011100101000110011001100110",
56 => "10100001101100011000101001010000",
57 => "01001100011100111110001000000111",
58 => "11010110001111100110001100001011",
59 => "10001000000001011010010111101010",
60 => "10011011101010010101110011100000",
61 => "00000110011111001000110011110101",
62 => "11101001111100011000110100010110",
63 => "01111111011100011011001011010110",
64 => "10101010100010010000000100110001",
65 => "11000011110011010011100011010100",
66 => "10100000111001111100010001010111",
67 => "10000010001110101110100011110001",
68 => "11110100000111110110000001001111",
69 => "00001010111111001101010011100100",
70 => "00110110111011110101101100110010",
71 => "01100101100011100101001001010010",
72 => "01010110011000101011011000000101",
73 => "11110101101011110110011101101011",
74 => "11001110111101101111010111101111",
75 => "01110101110101001000011001110010",
76 => "11101110011101001100101001111011",
77 => "00110000101111001100110010000101",
78 => "00111000010100011011111010100101",
79 => "00001000111101101000101000110011",
80 => "01000000111010000110000111100011",
81 => "11101010001110101100011110011010",
82 => "00010100101100010100110110011001",
83 => "10001001110000011010110001111111",
84 => "11011000000010001001100010111000",
85 => "10011010111101000100101100100101",
86 => "01000001111100111110111111000100",
87 => "10000001100100010000101010011110",
88 => "10111001000001100000111101000100",
89 => "00001010011100001110110000010111",
90 => "01000110010110111010001000010000",
91 => "01010110100110111000001111011011",
92 => "00010110000001001010100010100111",
93 => "01111000111100110110011011001110",
94 => "11010011000001111001011001101111",
95 => "00000001000010000011011010001010",
96 => "01101001010110001101011001110100",
97 => "10001010111011001100100011001100",
98 => "00111111101000100110010101101011",
99 => "00010100111100100010110000100000"),
(
0 => "0011000101110011001111101Y001000",
1 => "111101000000001110111101000010Y0",
2 => "000110Y1010100100101011111101011",
3 => "01100110111100101100010110000Y00",
4 => "01001001010110110110000111111Y00",
5 => "1010110Y101111101011010001000011",
6 => "1Y111000101011010010111001100111",
7 => "01001011110111001Y01111001010011",
8 => "1100011010011101010000Y001100111",
9 => "101101Y0001010101000010000001010",
10 => "001111100011011011100100010Y0011",
11 => "001001100Y0110010000001000000011",
12 => "0000000000Y011010101100000100111",
13 => "10111100001111100011Y10101111110",
14 => "0010101110Y100010111111100100110",
15 => "00000100111Y01000000110011011011",
16 => "0001111100000001Y000001111000000",
17 => "1111010101000001011111Y011010110",
18 => "001011000100011100100Y1110011011",
19 => "0111Y111111011101010110110110111",
20 => "001100101000111110010111111010Y1",
21 => "000110101110111Y1011001110110111",
22 => "1100100111010011010Y011001111101",
23 => "011010000010110101110111100000Y0",
24 => "01101000011101010011Y10011011100",
25 => "0001000100100110011110010100010Y",
26 => "01000Y10111000001100010010111000",
27 => "011000000Y0110010110010010000101",
28 => "01001110100111011001101Y00010111",
29 => "1111101000010Y010000011100001011",
30 => "10000001110Y10111010100110000101",
31 => "10110Y00011001011001001101000100",
32 => "011110010001011100110000010110Y1",
33 => "011101111001Y1011000000101110111",
34 => "001111011110111101011100010Y0100",
35 => "1001Y111101001000000111111100100",
36 => "1111001011111110011001011000010Y",
37 => "0011011010110Y100001001101000001",
38 => "0110001100Y001010001011101110110",
39 => "1000000110110000100Y010000101110",
40 => "00010111100100000001Y00101001010",
41 => "111001011111Y1110101011110111110",
42 => "0011111001010000101110010Y010001",
43 => "100000101000111110111011110011Y0",
44 => "00010000110000001Y10100001000011",
45 => "1011011Y110000111111111101101011",
46 => "100011101Y0100010010110111110100",
47 => "1111001Y000100100101111000101111",
48 => "0011101100001Y110100110111001100",
49 => "1010100011000100010Y000011111011",
50 => "110110001010110010010Y1011001111",
51 => "110100100111Y1111110000111101100",
52 => "1110101101100Y010001110100000100",
53 => "11100000011111111Y00001100110111",
54 => "01010100111011000010001111Y10100",
55 => "001010011000Y1100110001000000110",
56 => "10110100000101010100110Y11101101",
57 => "111100111100110011000011000Y1011",
58 => "0Y001110110110001110101111000000",
59 => "1000000110000101100010000Y100100",
60 => "1010011Y111010001100100000101101",
61 => "1101100011110000100010Y111100011",
62 => "01110000111101Y01101110110000111",
63 => "000001101011011110Y0111000100001",
64 => "11011000010111111100100110101Y11",
65 => "011111100011110100001001Y1000110",
66 => "0111110000100Y010011110110101000",
67 => "0111101110Y000000111100111011001",
68 => "0111101010100101000010Y001101001",
69 => "0101001100011Y011010011010111001",
70 => "010000000001000000000001001Y0000",
71 => "00011011Y11011111010111100010111",
72 => "11100Y11000001001110011010000010",
73 => "100001100111111000010Y0100000110",
74 => "000100001010Y1110100011010000101",
75 => "110000001111100Y1101111101011000",
76 => "001001101101101000011011111Y0010",
77 => "1011Y010101111110010110100001101",
78 => "00Y01111101101101010111000011000",
79 => "110101011100001111000110101Y0000",
80 => "1111000110011101001000Y101101011",
81 => "0110101101100001111001111001Y010",
82 => "0001011000001Y010111011010100001",
83 => "11111101001110001100100Y01001010",
84 => "01110011001111010Y10101100010011",
85 => "11010110010011100011Y00111111100",
86 => "010111110101011010000000Y0001111",
87 => "0011110111111111010011100011Y110",
88 => "111Y1011010101101111000000111111",
89 => "110101111010110010Y0001001000111",
others => "00000000000000000000000000000000"),
(
0 => "110111101010110110010110Y000Y011",
1 => "1101Y10110011011100011Y100010001",
2 => "010010111001000010110001101100Y1",
3 => "1111001Y0001Y0111011111100001010",
4 => "01100100111010100Y1011110101Y110",
5 => "0100Y0100100101010000Y0000111111",
6 => "1111101101010000Y1Y0011001100101",
7 => "101Y101001000101010Y100101010000",
8 => "1001Y00110110110111110011Y100100",
9 => "1001000110100Y00Y101000000000101",
10 => "1101001110101100011110Y1Y1101010",
11 => "1Y0100010000000000011000111Y1100",
12 => "00110101011110Y0Y100101010110011",
13 => "01Y01011Y11000000101100010000111",
14 => "000011Y10000101Y0010010010001101",
15 => "11011111Y100011110000000010Y0011",
16 => "001011000100110011000Y10Y1000000",
17 => "000YY010101001010011010001001001",
18 => "001110Y01Y1101110111100010110000",
19 => "00011000100010010Y000Y0111010110",
20 => "0011000010110101Y01100011Y011000",
21 => "01Y01011110110100Y11100010010001",
22 => "00001100010110101100YY1100001111",
23 => "0111001101000Y10Y011000110010100",
24 => "10000011101001011Y1110Y010011100",
25 => "11100111001000100111111100YY1110",
26 => "11010011000111100Y10100111000010",
27 => "011001100100100Y00000111010000Y0",
28 => "110011001100000000Y100000010111Y",
29 => "1010101Y1110100111Y0000000100100",
30 => "011111110000011Y01101010010111Y1",
31 => "00101100111011011111101Y11010Y11",
32 => "101111001Y0100000Y10110011100011",
33 => "00000YY1110110011001011011101001",
34 => "11101Y010000100010101Y1001011111",
35 => "00011100011010101Y010101100Y0111",
36 => "01101111111110101011011Y000010Y0",
37 => "100111111001101111110Y100Y010001",
38 => "100011000101Y1110100000110100Y11",
39 => "10111011110101110Y01010Y01100011",
40 => "01011010001Y0Y110010100110101110",
41 => "111111Y000000101101111010110100Y",
42 => "01Y0011111011111Y001000111111010",
43 => "000000Y010010000010101110001000Y",
44 => "0101010010000011111Y10100Y111100",
45 => "0111011Y0100Y0001100110000111000",
46 => "1Y000100110110001Y00110110000100",
47 => "111Y100101010001100110101011011Y",
48 => "111111111Y100Y001001011100010100",
49 => "100001Y0Y11101100101010100111100",
50 => "1101000101001Y11001Y101001011100",
51 => "11Y0111001000000101Y011010000101",
52 => "010010011111001000011110011Y1Y11",
53 => "1000111110011Y011100011110010100",
54 => "1Y01Y110011001100000100100111101",
55 => "000101000Y0Y11011010001010010100",
56 => "10Y10100110Y01110101110010001101",
57 => "110Y1111111100111010Y10001101001",
58 => "11000011Y01001101101100101Y11100",
59 => "01011011100000101010Y0111Y000111",
60 => "00101Y101Y0001001011011010000011",
61 => "01101010111101110Y0000111101Y000",
62 => "1101000101010Y01100100101101Y111",
63 => "10101Y00101110111111Y00011110111",
64 => "0011010Y101111101010110001Y00111",
65 => "100100YY111011110111000101000000",
66 => "1010100Y010110100010001000101001",
67 => "100110111100111011101011Y000111Y",
68 => "00100Y00010000011Y11101111011000",
69 => "11100000010100010100010Y01000Y11",
70 => "00Y111101111100110Y1110110011010",
71 => "1Y11001000001000000010111110001Y",
72 => "1000100101Y111000111101Y01110110",
73 => "1111111010111Y1000Y1011100110110",
74 => "00010001Y010101000011Y1101000110",
75 => "1100Y000001000111101Y01001000011",
76 => "000011101100000000111Y1101101100",
77 => "0010100Y100010011111111000Y01000",
78 => "100010110110110011000101111Y00Y0",
79 => "00110011111100101111011YY0011111",
others => "00000000000000000000000000000000"),
(
0 => "011011Y001010010100111Y0Y0010000",
1 => "01100001100Y1011111Y0Y0100110111",
2 => "1001011110000110011011Y1110001YY",
3 => "10Y011011101001Y1001111100Y11110",
4 => "011100Y1011111010Y0110100111100Y",
5 => "1010Y00000000010111110110011YY10",
6 => "1Y01Y00000Y111110011100001010001",
7 => "0110Y1101100101001101Y1Y11101010",
8 => "00011Y00Y001100Y0000101000100010",
9 => "0010110110001010Y011Y1000Y101101",
10 => "1Y1010100Y11000Y0000000101001010",
11 => "011100Y00Y000010Y111111111010100",
12 => "0101001000110Y00100Y10011111101Y",
13 => "110011110111Y011110Y0101100Y1100",
14 => "1Y01001100011Y000011Y10100011110",
15 => "0111101001Y0100Y10000100101Y0000",
16 => "011111110100Y110100100101Y110Y10",
17 => "1010111010000000010100001111YYY1",
18 => "010000110011000001Y0Y001Y1110010",
19 => "1011110001Y0YY110000000111100101",
20 => "110111Y0010110Y0Y000111101010011",
21 => "01Y010001011010110110Y1110111Y00",
22 => "000000Y01011001Y0010111111Y11011",
23 => "01Y00000100Y001011Y1110001001100",
24 => "11001100Y01011010Y01100101110100",
25 => "11100111011111101Y1111010000YY11",
26 => "001010101Y100101111011Y100011Y01",
27 => "01Y0101100Y1111000100000Y0001101",
28 => "0Y010100010100010Y0Y111010110111",
29 => "1000011111010001Y00Y0011111Y1011",
30 => "101011111001001Y00Y0Y00101101000",
31 => "10101Y00000000111100Y111Y1101111",
32 => "01001000Y10Y1101101Y010111101110",
33 => "0110001100110100011011Y0Y1Y00011",
34 => "10101Y0000100001111Y111001111011",
35 => "01001100011001100Y00Y0Y001100001",
36 => "1110010110111Y0101001100YY100110",
37 => "1000001010YY0001101100001000001Y",
38 => "011010000100Y000001000Y10Y100010",
39 => "000Y111010100100Y1011Y0111111000",
40 => "000010000Y00Y10011100Y1011100110",
41 => "1100111011001001111010010Y0001YY",
42 => "0110101Y1001100111011Y000000Y111",
43 => "101100Y0100101110Y1011Y000110110",
44 => "1101Y111110Y0001001Y011100011001",
45 => "01Y0Y101011000100111100111000010",
46 => "000011100Y101Y000Y01101010100011",
47 => "1Y1110111110Y11110100000100Y1001",
48 => "0000100Y01100000110100Y010001Y00",
49 => "010Y11000100100011100Y101111011Y",
50 => "0100Y11111101000010110Y001011001",
51 => "1Y1Y110011Y011110010100011111101",
52 => "01101011Y1010Y10010Y000001001001",
53 => "1Y00Y10010001100100001111Y111111",
54 => "000Y111110110Y101010001Y01110011",
55 => "01111Y110010001010101YY000011111",
56 => "01000000111Y0000010Y00001Y100101",
57 => "100110Y111110100Y11000Y000111011",
58 => "0101100011111Y01110001Y1000010Y0",
59 => "0000010Y1000100110100YY010111000",
60 => "1111000100100000001YY1Y101101110",
61 => "110000Y0100Y100000111001100Y1100",
62 => "00101001010100001000Y1001YY01010",
63 => "0000101Y100101011Y110010Y1001110",
64 => "1Y00100000010Y010001110001Y00010",
65 => "11010Y10001100Y01001000000100Y11",
66 => "10010101101Y0101101Y1100Y0110111",
67 => "101Y10011Y0101101011100100Y01110",
68 => "0Y110010001110Y0001110Y110011101",
69 => "1011001Y011Y1Y010001101100101011",
others => "00000000000000000000000000000000"),
(
0 => "101000000Y1110010Y01110110YY1111",
1 => "1100110Y1000010Y111001001Y00100Y",
2 => "01100Y11000001000Y0Y010Y00100010",
3 => "0Y001000010001010110110Y100Y010Y",
4 => "0101100111110Y0101Y1Y1011100Y110",
5 => "010Y0Y000000111101010Y0Y11110101",
6 => "010110Y0Y0100100010101000Y101011",
7 => "011101100Y0Y11110011000YY1111111",
8 => "11Y110Y1Y1100111Y100001101110100",
9 => "000100YY011Y110100101101111110Y1",
10 => "01101Y1001Y00000000010110Y00Y101",
11 => "10Y11000110Y01011000010000Y000Y0",
12 => "10Y01Y00001111101Y111110000Y1100",
13 => "11011100110000111Y0001000Y1Y10Y1",
14 => "0101100011Y000YY111110100Y100001",
15 => "101111100Y00001Y11Y101110Y110110",
16 => "1111111111101011100Y010Y1110Y100",
17 => "11101110Y000YY110001110Y11000101",
18 => "010Y0100110Y01001Y1011001100Y110",
19 => "110000001100Y11Y000Y1011Y1101011",
20 => "1Y1010001YY101010Y11100110011110",
21 => "1101011011101Y00Y101000Y00101Y10",
22 => "11Y00Y100Y0011Y11101111011101011",
23 => "1101000101010010101000YY100Y1Y10",
24 => "101Y001001100Y001Y11Y00110011000",
25 => "11Y101100Y01110Y0101001000100Y01",
26 => "10101101Y01110110Y0Y00111Y100001",
27 => "011111Y01111001111Y110Y010111Y11",
28 => "0101100Y1Y10011011111111YY010000",
29 => "00001Y101111Y1Y11Y10100001010111",
30 => "110Y0Y100Y10000000011111110110Y0",
31 => "00100Y10011Y0000001111Y1Y0010010",
32 => "0101010Y1010000011100Y0110101Y10",
33 => "110000YY10111101101001001Y0Y1010",
34 => "110001111Y0001Y001101YY000000011",
35 => "001Y0100011011Y0Y0Y1111110110011",
36 => "1111011010010101Y1YY0111Y1111011",
37 => "1YY11101010000Y1010110001010Y100",
38 => "001001YY00011110000100111000Y100",
39 => "01110000001101Y1Y01110Y0011001Y1",
40 => "0101Y00011Y01111101110Y111111101",
41 => "1Y10Y0Y110110000Y000110011110111",
42 => "001001Y1111101Y1101Y111100010Y00",
43 => "1Y00Y0100101010001100Y0001Y00100",
44 => "000111Y01100010001100YY100001Y00",
45 => "1101Y11Y010Y11Y11000001111010100",
46 => "01000000001Y1YY10001110110Y11001",
47 => "0110101101011Y1Y111Y111100111Y11",
48 => "01010110011001010001Y10000YY1011",
49 => "00Y1011Y1101011100Y01010001111Y1",
50 => "0Y1011Y101100010Y0010100010Y0101",
51 => "111000Y0011011110101101Y0010Y00Y",
52 => "1Y01100010001Y1001111Y11100100Y0",
53 => "0Y01Y01Y0Y1011111110011110010101",
54 => "1Y00Y1Y101001000001001001011101Y",
55 => "100111Y1010001001100101YY0Y11010",
56 => "000Y1111111100Y00010Y110011Y1101",
57 => "1111100101Y001Y110111Y0010000Y11",
58 => "000001010Y100010000001Y00Y000000",
59 => "010Y01Y10100010110111Y111010Y111",
others => "00000000000000000000000000000000"),
(
0 => "0011111000Y1011Y001Y000111YY0111",
1 => "01YY000011Y1101100001Y110110Y110",
2 => "01Y11Y1111Y1000100000100Y00101Y1",
3 => "1011Y001Y1010000111Y10011Y0Y0011",
4 => "0001110Y011010Y00YY110101110111Y",
5 => "000YY101YY1100110010110111101Y11",
6 => "1101111Y101010Y111001Y0111001YY0",
7 => "1000100101000Y10YY1100Y101011101",
8 => "10111Y0110001Y110Y011Y1001Y11110",
9 => "1001101110Y010Y1100Y10001111Y001",
10 => "011111Y00111Y011Y111100YY0100010",
11 => "0101Y1100010001000001Y0Y1YY10001",
12 => "0011110Y1100Y0011111YY100Y100010",
13 => "0010010Y00110000Y0001111Y1101Y1Y",
14 => "1010001001010YY01Y110Y001110Y001",
15 => "1Y0010111Y1000110Y10Y001010100Y0",
16 => "010011Y1011001001101Y0YY0110Y101",
17 => "01001Y001000101000YY0Y1101000001",
18 => "011100011Y001Y1000110Y0010000YY0",
19 => "00111Y0011001001Y11Y011110YY0100",
20 => "1010001110Y011Y001Y00011Y10101Y0",
21 => "01000101Y10001Y10Y011111Y0110001",
22 => "0100101Y01Y000001010Y0Y00100Y001",
23 => "0011111YY101Y0111011101101110100",
24 => "01001011111Y0Y1000100011Y011111Y",
25 => "0011110Y01110YY0010100100Y100000",
26 => "0100111Y001Y1Y101Y11001100101001",
27 => "10000Y11001Y11Y00111111101Y01111",
28 => "101100YY1Y01011010Y1101010000100",
29 => "0100Y100Y0100Y0Y1Y00000001010011",
30 => "00Y011000101Y100001101Y101100Y1Y",
31 => "1100100Y00Y0010110Y1110Y0011Y001",
32 => "0Y1Y0110000Y1111Y1000011111011Y0",
33 => "0100110Y001Y1000Y101001001Y10010",
34 => "1110Y00YY1101Y10011010001001Y010",
35 => "0011001101001000Y0Y1Y110Y110001Y",
36 => "001100Y0010110Y110100101Y00Y0Y01",
37 => "01000000000010001000Y0YY100Y10Y0",
38 => "1Y1101Y101110Y101010011100Y10Y00",
39 => "1000Y0Y1110Y011000010Y0001Y10010",
40 => "11YY0010011110Y0110Y101111000Y01",
41 => "110111101010010Y1Y1YY0Y111100010",
42 => "0001Y011110Y000YY01Y110101010110",
43 => "01YY0110111Y00011Y1001111100Y111",
44 => "1001Y0001100Y0YY11101Y1001101001",
45 => "110000100001110101YY010101YY1010",
46 => "1000111Y000000111Y101Y101Y1000Y0",
47 => "000YY1Y000000110000Y10101Y110100",
48 => "100101000Y001Y1100100Y01101Y000Y",
49 => "111Y1010011Y1010YY10101111010000",
others => "00000000000000000000000000000000"),
(
0 => "0Y10000110Y101000110100100Y10Y1Y",
1 => "011000Y10011YY000Y000Y01Y1011111",
2 => "00001011010Y0YY0111Y10001111Y10Y",
3 => "101110001110101Y0YY11000010111YY",
4 => "110101011YY10Y01Y11001001Y000Y10",
5 => "00Y0110011011010100Y001Y1001YYY1",
6 => "01Y11110Y0Y1001100101Y1Y0Y111010",
7 => "1000Y11010011010Y1010YY00YY11100",
8 => "001010YY1Y1111Y00011001000111Y0Y",
9 => "1010011001110YYY1100000Y10111Y11",
10 => "000Y1100Y10001Y111010101Y101Y00Y",
11 => "11Y10011Y0101110Y0Y110Y0111Y0110",
12 => "11100Y1YY0111YYY0001000101000111",
13 => "10101Y000100Y11Y01Y1011101Y010Y0",
14 => "101011010Y101Y10Y00Y10100Y100Y00",
15 => "111YY010111100Y11Y010000Y1Y00101",
16 => "01110Y0011Y1010Y111Y1010Y0011101",
17 => "101000011YYY1011101Y10001Y1111Y0",
18 => "11101Y0001Y1Y001011001Y110Y100Y0",
19 => "1Y1111001Y1101Y001Y1011Y11001101",
20 => "011Y101Y00101Y111110YY0Y01000110",
21 => "110101010YY100011010100000Y1Y001",
22 => "10110100101Y110Y11011Y0Y0YY10001",
23 => "011100101111Y100YYY0111000Y0Y001",
24 => "01Y0100Y1100Y000010Y10101Y010Y11",
25 => "011Y1010Y0Y0Y00011010000111Y100Y",
26 => "10001Y011011Y0Y01100Y0101001Y111",
27 => "0YY101010101101Y000Y1100Y1Y01111",
28 => "010Y01011Y00Y0100011011Y01100YY1",
29 => "0010001110Y0110100100Y01Y0YY11Y1",
30 => "010010YY00Y1000Y1Y10100011110Y00",
31 => "11000100010Y1YY0011001Y0Y10011Y0",
32 => "11110101Y1Y011100YY0110Y00Y01110",
33 => "0Y010010100010100Y11Y111011YY01Y",
34 => "11011Y1000110111Y10101Y11011Y101",
35 => "01Y0011010Y001100000YY111100YY10",
36 => "01111Y00011Y0011YYY0011000010101",
37 => "01101010Y0011Y100Y10000YYY111011",
38 => "0111Y0YY0Y111Y010010100111101001",
39 => "1101010Y00001111101YYY1Y100Y1011",
others => "00000000000000000000000000000000"),
(
0 => "1YY1000100110Y110YY0YY0100011100",
1 => "1Y1101001001001Y00111YY0Y0Y10011",
2 => "110Y0YY0010101Y001101Y111101000Y",
3 => "11Y001101011Y10Y11Y011YY11010101",
4 => "110Y111Y1Y00001101Y11111001YYY00",
5 => "10Y1110YY11010YY0001Y0Y110010101",
6 => "11Y111Y1110101110101Y10100YY001Y",
7 => "11Y1000Y111Y100010001YY11011Y00Y",
8 => "10Y0011Y0110Y00110Y0100Y10Y000Y0",
9 => "1000101011Y10Y11Y110Y01Y1YY01011",
10 => "00100Y1Y1Y0110Y10100010Y10010001",
11 => "1Y100110Y1000Y0Y100Y001101Y00001",
12 => "0000100Y1000YY000Y0001Y00110Y00Y",
13 => "101100Y110YY10001100YY011001Y000",
14 => "110Y10000110Y00Y101101Y00100011Y",
15 => "11100Y11YY101100Y0Y100001Y0011Y1",
16 => "01000Y1Y011000Y10101Y1110YY0Y011",
17 => "1Y010YY11101101Y10Y10Y0000100001",
18 => "111Y1Y00110110YY00Y011YY10111111",
19 => "00111Y01110Y1011001110Y1100YY1YY",
20 => "11111Y10Y01011000011Y00Y01Y00YY1",
21 => "100Y111101YY00000011Y001Y0Y11001",
22 => "0YY0000Y110101100000Y10011Y111Y0",
23 => "0Y01000Y01100100100Y11111Y101YY0",
24 => "1100Y1111000011010Y0Y1001Y0YY0Y0",
25 => "00YY11111Y10Y0100011010010Y1Y010",
26 => "0Y000100Y100Y001010011011Y1Y0Y10",
27 => "1Y101100YY0Y0100Y011100010100YY0",
28 => "001Y0Y110101Y01101001011001Y01Y1",
29 => "0000Y00YY1100000011YY10001Y1111Y",
others => "00000000000000000000000000000000"),
(
0 => "0Y10YY0111001010Y1Y0010101101010",
1 => "1001011Y1YYY11000Y0111010011YY0Y",
2 => "10011Y01Y1110Y0111Y10Y10Y010YY11",
3 => "1Y0011Y00Y0Y00Y0001110Y011101001",
4 => "0Y011001010Y1Y110011Y01Y10001Y01",
5 => "10YY111Y011Y1Y0111110Y1110100Y01",
6 => "010001Y1Y1010Y0YYY1Y010001110111",
7 => "000Y1Y00Y11111000111Y10YY100Y11Y",
8 => "0100YYY1Y001001111Y11Y01010Y1101",
9 => "0010001Y11001110Y10Y0Y111111Y0YY",
10 => "0Y0000Y1010Y0Y010101YY1110001100",
11 => "1Y011Y010Y10111Y0Y10Y11110YY0100",
12 => "01Y11010Y1000Y010Y0100110010Y0Y1",
13 => "0Y011Y110Y101011011Y100011Y0Y001",
14 => "11000010Y1Y11YY1Y0Y001000YY10000",
15 => "1001Y0001YY11Y010Y11Y1Y000101Y10",
16 => "00000YYY1101100Y0Y11YY10000Y0111",
17 => "0000011Y1101001Y0YY1010YYY011000",
18 => "11YY1101YY0Y1110101000010001Y111",
19 => "0Y10110010Y0YY000001000YY0Y0011Y",
others => "00000000000000000000000000000000"),
(
0 => "000Y0001Y010Y1YY1Y1YY000Y0011101",
1 => "111Y10Y1110111YY0010001Y010Y1YY1",
2 => "010Y0110Y1110YY11YY1110110000110",
3 => "01Y111Y1111Y11Y11Y1Y000Y111YY000",
4 => "1Y11Y10YY0Y10Y10Y10111YY11100011",
5 => "10Y01YY1100111010Y111YY01Y01101Y",
6 => "011110111Y01010YY0YYY11100Y1YY00",
7 => "00Y1Y11Y1100000Y01Y01Y0111Y10001",
8 => "01Y101Y0Y111Y11Y0100101Y001YY001",
9 => "0Y0Y1Y0011Y011Y1Y1Y110111Y10Y010",
others => "00000000000000000000000000000000"));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;