library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => "01101111111110111111111111101011",
1 => "10001110111011100110000100101001",
2 => "10011010001010111001111011000011",
3 => "10010011010101100001101011000010",
4 => "11010100111110100000111011100100",
5 => "10100101100010110101000111111110",
6 => "00111111011110001010111101110010",
7 => "10001001011100100000101011100111",
8 => "11010111010001000000101110101110",
9 => "00101111101010001011001100001101",
others => "00000000000000000000000000000000"),
(
0 => "000101010100110110100010011010Y1",
1 => "011110011010111110001111111001Y0",
2 => "00001110100111101Y11000100010101",
3 => "00110110010Y11011001101100001000",
4 => "00011110110Y11000001011110110011",
5 => "0010111110111010Y000100000100010",
6 => "00010110Y11100100000011001110110",
7 => "111011011001Y1100111010110010101",
8 => "10000Y01011110100101111001101100",
9 => "01101011100100Y10111010111000101",
others => "00000000000000000000000000000000"),
(
0 => "1100111Y101001101100Y11111100100",
1 => "111Y110011101101011001110000001Y",
2 => "111101100101001Y100Y011101010011",
3 => "01000Y1010Y011110100100111001011",
4 => "1011Y01111101Y010010010000001000",
5 => "1110000110100101101Y1110100110Y1",
6 => "0010011111111010001Y00111000Y001",
7 => "1Y000Y00101001111010010101101110",
8 => "000111110Y11000011101011110Y1011",
9 => "110110Y010110010110000000110Y101",
others => "00000000000000000000000000000000"),
(
0 => "1000101011010000Y1Y11000Y1001100",
1 => "1101010010001111YY011110000010Y1",
2 => "01Y11010101001101111Y1101Y011010",
3 => "010111010000Y01101111Y000110Y011",
4 => "0010101Y0011011Y001Y000001011100",
5 => "00011100000Y00111101Y01Y00101111",
6 => "01001001011Y100001Y1110Y00011110",
7 => "010000Y00110011101000000Y111Y101",
8 => "010100100110000010000Y110000011Y",
9 => "0110010100001Y11100000100YY10000",
others => "00000000000000000000000000000000"),
(
0 => "101Y1010Y1Y01111000001Y101110010",
1 => "11011010100Y1Y0100101Y1001001110",
2 => "01011001100Y01Y1111Y11101011Y011",
3 => "000YY11Y11110110000Y111110111100",
4 => "0111Y010Y10101110010YY1011001111",
5 => "01111001101100Y10110101Y0Y01Y010",
6 => "0Y111110011YY0111Y10011111110011",
7 => "1Y11001110Y011001Y0100001011Y100",
8 => "01011000Y00011110100Y011010Y111Y",
9 => "100Y10Y0Y10011001100010011110000",
others => "00000000000000000000000000000000"),
(
0 => "110Y01000010010111Y1111110000Y1Y",
1 => "111111010110Y11Y0Y10110011101YY1",
2 => "01Y00Y10Y11Y11Y10111000110001011",
3 => "0010001111Y0Y000111Y110010Y10011",
4 => "101010Y0Y010001000111001Y0Y10101",
5 => "0100000YY0111101Y0Y0101Y00100110",
6 => "10100010Y0100YY00100Y11000111100",
7 => "10Y10Y01100YY11001001010Y0110101",
8 => "01110001Y000000101Y11YY11101010Y",
9 => "1101Y00000111110001110111YY10Y00",
10 => "110Y01Y101Y110010110Y11111111001",
11 => "11100101Y00100Y01Y10000001Y00001",
12 => "111YY100Y11001Y011110Y1010010111",
13 => "100Y0110Y11000100Y0Y100011000101",
14 => "10100Y01010100111Y0110100Y11Y1Y0",
15 => "00Y1011011YY001Y0111000001100101",
16 => "00Y10110000111Y1011Y0Y1101100111",
17 => "01Y0Y10Y010100110101011101010Y11",
18 => "110Y001101YY000010110000Y1111010",
19 => "0Y00001100101001000110011Y1Y1YY1",
20 => "1111Y00010101000001011Y010Y1Y010",
21 => "00000Y111001Y10101Y1101YY1001010",
22 => "11001000010Y10010010Y0010Y1Y1101",
23 => "1Y111110Y10101011YY011100100011Y",
24 => "100010001000Y10111Y0Y10Y1001Y101",
25 => "101101010111Y10Y0Y110111100YY111",
26 => "00Y0001Y00101011101100111Y01111Y",
27 => "0001011010Y1111101Y0Y0100011Y0Y1",
28 => "001110Y010Y111011Y1110Y111111Y01",
29 => "011001001Y1YY0110100000Y00Y00000",
30 => "11Y110Y0111111Y1Y111011110Y10000",
31 => "001011111Y1Y01111Y10Y101000101Y1",
32 => "10Y01000Y000Y10101001001Y0Y10000",
33 => "010011101110Y101101Y0Y1000000Y1Y",
34 => "0000110Y001Y111Y01Y1001Y11001010",
35 => "110Y1YY11Y0111101010111110110Y00",
36 => "100Y0Y0Y0010010Y01000010Y1100111",
37 => "1010Y10000011Y11Y00010101Y1Y0011",
38 => "1001011Y00010100Y100011101Y1Y1Y1",
39 => "0Y0011YY011YY1001010101100101000",
40 => "1110Y001011111011000Y00Y1Y010Y11",
41 => "001Y01YY110Y1101Y110110001110011",
42 => "0Y011Y11Y001Y1110110111011Y00111",
43 => "0Y00011Y1000011YY00000000110Y101",
44 => "0011000110Y101Y0Y00Y1010100101Y1",
45 => "0011Y0100010Y00Y000YY10111000011",
46 => "10Y001Y0010101Y001Y111Y001010010",
47 => "0YY000100111Y1010100100111111YY0",
48 => "11Y11Y111Y1Y1Y111011101100100100",
49 => "111YYY000011001Y1010111110Y11010",
50 => "0Y01101111100110111YY1001001Y010",
51 => "111YYY010010Y0001001010Y01100010",
52 => "110Y0111011100Y1111Y01110111Y001",
53 => "10111Y010011001101Y01Y101Y10111Y",
54 => "001101101Y0Y0011Y001000001Y11Y10",
55 => "11Y01110101Y10000YY1011100011100",
56 => "11001010010100Y1110011Y1Y1111YY1",
57 => "010Y001100Y011010110Y01Y0011Y001",
58 => "010000Y1Y01Y1111Y00010010100Y101",
59 => "101101Y01Y0000011111001Y0Y0Y0001",
60 => "100Y0011Y001101Y1000101011YY1111",
61 => "11011Y01000Y00Y1Y01000100011Y100",
62 => "10Y0Y0001011001Y1111100010000YY1",
63 => "10100101YY10Y011000Y1000Y1001111",
64 => "101Y110001010110Y0Y00Y11Y0110100",
65 => "0Y011001000000Y10101Y11001011YY1",
66 => "101Y10Y1001111001Y000011110Y1001",
67 => "0010011001101100010100Y10110Y0Y1",
68 => "111100Y11111101100Y00111Y00Y00Y1",
69 => "10011010101Y00110Y0101YY10001110",
70 => "001Y10110100001011YY01010Y0Y1111",
71 => "11YYY100Y10101011100011101111100",
72 => "00YY001101111Y01010011Y000111101",
73 => "1Y11110110Y01010Y110001010Y11011",
74 => "11110010000Y100Y0110Y101001Y0100",
75 => "11111000110001010Y11YY0010Y10Y11",
76 => "00000101010Y0Y1Y1010111100Y1010Y",
77 => "1001110100000010Y10Y1100Y100100Y",
78 => "1010110YY01101111011Y01011YY1100",
79 => "00111010001110Y11001100YY010100Y",
80 => "11Y1Y110Y11000Y11010Y11111111101",
81 => "0Y0110Y001101001Y0010Y10Y0100111",
82 => "1000100100Y01011Y00Y00101YY01101",
83 => "10Y110010Y1Y11Y0Y110010011111110",
84 => "0Y1YY011000001110Y01001110000Y01",
85 => "0100101Y0Y110000YY1Y100111111110",
86 => "110Y10Y10010000100Y01Y1Y00101010",
87 => "00000Y1Y0Y1111110Y0Y100011100100",
88 => "10101100011000101YY111YYY0100100",
89 => "00Y11001011100001Y001Y11Y1110001",
90 => "0Y1001111011001110011Y1111YY1101",
91 => "010Y0Y000011010Y000001100Y0101Y1",
92 => "1Y101111100110Y100Y0Y1Y100000010",
93 => "10Y0Y11Y1Y0010001110010110011Y01",
94 => "101001Y10001YY0110000110001Y0111",
95 => "000011100010Y01YY11011Y111Y01011",
96 => "00Y01Y0110010100100000Y00Y110101",
97 => "1111Y10Y01Y010010111111001Y0Y000",
98 => "111Y11Y010000000010Y0Y111Y110101",
99 => "1Y101110110111Y1101111YY0Y100111"),
(
0 => "00000111110010YY100Y0010110Y00Y0",
1 => "10110100YY1101Y111110Y1011110Y0Y",
2 => "0001Y11011Y111Y000110101YYY01100",
3 => "01YY011101001Y01011Y000010YY1110",
4 => "010110000010Y01101000YY00Y1100Y0",
5 => "01Y1Y010100Y111YY110Y11101101111",
6 => "001101Y0110110YY1110101YY10001Y1",
7 => "01000111Y1Y00110101Y1111Y10111Y1",
8 => "101Y01001100010Y0Y010Y0Y01001Y11",
9 => "01Y1100YY1011111101Y0111011Y1101",
others => "00000000000000000000000000000000"),
(
0 => "010Y1Y1Y0Y011Y00011011Y111010101",
1 => "10101YY0110011001Y000Y001100YYY1",
2 => "001001001Y0Y1001Y10Y000111YY10Y1",
3 => "11100101111Y1Y010Y1Y110Y110100Y1",
4 => "10YY100111Y1001011101010Y1YY0100",
5 => "11011Y00Y0111100Y1YY0111011101YY",
6 => "0001111101Y1Y010111Y01Y11100Y0Y0",
7 => "1Y10Y0011001Y0110Y110Y110Y10Y000",
8 => "01011110Y11Y1YY011000Y00Y011111Y",
9 => "00YY001110Y01000Y0111Y1Y1001Y111",
others => "00000000000000000000000000000000"),
(
0 => "1Y011Y0101101Y10Y1111Y1Y100000Y0",
1 => "0001101Y010101Y1Y1000Y01Y010Y00Y",
2 => "1Y11000111011YY1Y011Y00Y11Y0010Y",
3 => "0Y0111YY11Y111Y11Y1Y0Y1111111100",
4 => "00YY101Y1011110Y011YY111Y0101011",
5 => "00Y1101Y0010000YY11111101Y00010Y",
6 => "0001Y10100100Y1YY100Y11011Y10001",
7 => "11Y1110Y10011Y0Y1Y01101Y101Y1001",
8 => "011YY10Y10Y110011100Y11YY01010Y0",
9 => "00Y1YYY00011Y1011Y01Y0100010110Y",
others => "00000000000000000000000000000000"),
(
0 => "10110110001YYY100000Y0Y1Y10Y10YY",
1 => "1110Y000000YYY10Y01111111101Y00Y",
2 => "0YY0Y100110110011110YY00Y100Y0Y1",
3 => "1Y01110Y1010111YY1Y1YY11Y0010010",
4 => "0101Y10110000Y0111Y110YY1YY0Y001",
5 => "101YY101101YYY111110YY1000001011",
6 => "1Y0Y00001111Y1000011YY100YY11100",
7 => "00000YY1010001Y1Y1111Y1Y01001101",
8 => "1Y001Y0Y1Y1110YY0011Y01Y10Y10011",
9 => "0Y1Y10100011Y1Y1YY0001010010Y01Y",
others => "00000000000000000000000000000000"));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;