library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM : TCAM_ARRAY_3D :=
(
(
0 => "10011100001010000101010110101011",
1 => "11001001010110010100110111100101",
2 => "10000101000011011010000110101101",
3 => "00110110100111101010111011101011",
4 => "00101010010111100010101111111111",
5 => "00111011001110000110001010101111",
6 => "10011110101101001111100000100111",
7 => "00111110001011010000100010110010",
8 => "10100100100000100101111001110100",
9 => "10111110010101000110111001000011",
10 => "01001011110010101011110111100100",
11 => "00000101101000010000100101100110",
12 => "01100000110111111010110000111111",
13 => "11100011011000100011111110010110",
14 => "10010110110111110100100010110011",
15 => "11100101110011101010110000100010",
16 => "11110000101011101010010101001101",
17 => "00101000100000000111001101001011",
18 => "01110010001101101010011111001101",
19 => "00001011100000010110001001101100",
20 => "10100100011001111001001000101111",
21 => "11011101010011011001010001111001",
22 => "00100100011011111001000101000011",
23 => "01111101011111000011100011101110",
24 => "11101110011000111100000101110111",
25 => "11010011101110100101001110111100",
26 => "11010010111111111100011010101101",
27 => "01110011010011111110011011011000",
28 => "00000010111001110111010110111101",
29 => "10011110110111111110100100101110",
30 => "00000110101111100000101001000010",
31 => "11101110000010010111000011111000",
32 => "00100110101001100001111100010001",
33 => "10101100001110001100001101111000",
34 => "00011101010010111011101100011011",
35 => "10010110011111101110000111111010",
36 => "11100101001000011100111101111100",
37 => "11100001011001000111111011110110",
38 => "00001110010010101111110000111011",
39 => "01011010001111001011111111110100",
40 => "10001111111100011001111011001010",
41 => "01000110011010010000110101111110",
42 => "01100010110101000110111101101000",
43 => "11000001010011111110001111010011",
44 => "01100010000000110111000010001000",
45 => "11010111111001001100000000110000",
46 => "01101011001101111011010111011001",
47 => "11011011011001111101111010011110",
48 => "00110110101011101100011111001100",
49 => "10100000000001111010111001100111",
50 => "10101011100010011001001000010010",
51 => "10010011001000111010000100001101",
52 => "01001010100110110001111110000111",
53 => "10011000101001100100101110001101",
54 => "00011010000110110011011011110111",
55 => "01110000110000100001011001011011",
56 => "01110110101100110111001000000000",
57 => "01010001100101000010110010000100",
58 => "00000000001101001110110100101100",
59 => "01011010001100100111100011001011",
60 => "11001010100100010110000100010111",
61 => "10000010110100010011000101011100",
62 => "10001111100001000100100100001010",
63 => "01100001000010010111111110010001",
64 => "01110100000111101100111010111110",
65 => "01110101100011010001001011011000",
66 => "10100000011011001100010011111001",
67 => "00101111100110111010110100000000",
68 => "10011011110010111011011110000001",
69 => "00100001110000101001010110110010",
70 => "00001011011010101011010000010011",
71 => "00011111011000011011001101000101",
72 => "11010000000011011111001000110010",
73 => "11001010000101110011010110101000",
74 => "01111000101100011111111010001001",
75 => "01100010001100101000100111010100",
76 => "10010011101000011111010001000010",
77 => "00011101010100100100111010010101",
78 => "11100110000010100000001001111100",
79 => "01110100100000101000100011110110",
80 => "01011100001111001110010011110111",
81 => "01010101000011100000010101110100",
82 => "10001001110000110100100111101001",
83 => "10011010101101010000101111110000",
84 => "11100110011101010010110001101101",
85 => "10001000000011010001111001110110",
86 => "10010010000001100000011111001110",
87 => "10010110101110000001000000111011",
88 => "01110000000110010010011001111001",
89 => "01110000010111000111000110111000",
90 => "01010001111010010101010110110110",
91 => "01001010001111001001001000011100",
92 => "11011111110011010010100110010011",
93 => "00100001101110110111010010001101",
94 => "11000000001010100000111100001100",
95 => "01101100010011010011111010101101",
96 => "10000101110101101100010011111001",
97 => "10001111111110111001111101010100",
98 => "00010101010010011111011111010011",
99 => "01110101110000000011101111100000"),
(
0 => "11000110001110010011101Y11000000",
1 => "10010100Y10110101101111011000110",
2 => "01111Y00000001110011000001011010",
3 => "011101010111011000100011010111Y0",
4 => "01111101110000101Y00001010111001",
5 => "1011Y101001111110101001100111100",
6 => "1100100111001101111001110Y001101",
7 => "0Y110110000010100011010001010010",
8 => "1010011010111010Y101110100010000",
9 => "11Y01001011011010000111100000101",
10 => "000100100011100000101000100Y1010",
11 => "01110010101111101111101100Y00101",
12 => "0Y101000111000100110101000110100",
13 => "0100011001001001111100000Y110011",
14 => "010111001111101000101010Y0100101",
15 => "000111110010111001001Y0000110001",
16 => "111101101Y0010001011100100010111",
17 => "0100111100011001001011011101Y000",
18 => "011101000011Y0000011111101101011",
19 => "00100110101010011000001Y01001111",
20 => "1001111011001000Y100001110000101",
21 => "00010111010100100110Y11010101111",
22 => "01101111010001101001Y11001011011",
23 => "0101001101100110000Y010111100001",
24 => "10011010101100110100111100Y10000",
25 => "00100110110011111000000101111Y11",
26 => "0110Y000110100101101110010001000",
27 => "011111Y1001000001111001010101110",
28 => "01011001Y10000110110111111101010",
29 => "1Y011101000000101000001111100111",
30 => "11010Y01000000101001001000100110",
31 => "0110000001110Y011111100100110000",
32 => "010111001001Y1001101010110101010",
33 => "1011011001000111110100Y010111101",
34 => "01101011Y10010110000100101111110",
35 => "00010Y00000010110001010001001110",
36 => "000100011000110110Y1100000111100",
37 => "00100010010111Y10101010001111011",
38 => "01Y11010110001110001001000001111",
39 => "10010001111Y01101100101101010000",
40 => "0110101001000000Y101000011001110",
41 => "0111Y100111010000011010101110010",
42 => "0100001100110Y001101111000001100",
43 => "00111100101011111001001011010Y01",
44 => "0000Y110010100110101111000111101",
45 => "10100111111011100Y10110100010001",
46 => "10010100000110Y00110110000110110",
47 => "00000000101100Y00011101010011110",
48 => "00000111Y00011101011110001110110",
49 => "01010100011111110Y11000000111110",
50 => "1000101110101011101001111010Y001",
51 => "010111110111001010011011010101Y1",
52 => "1Y000000110101000101110011110011",
53 => "00101010010010100Y10111001101101",
54 => "10000110100000011011100110110Y01",
55 => "000111010100Y1101000001100101110",
56 => "0101101011110001110001010Y101101",
57 => "1001011Y001110000010001001001011",
58 => "111Y1110100100110010100001010100",
59 => "10000001001101110000Y00101111010",
60 => "1011111Y100001000010100100011010",
61 => "10111111110011111101001001Y00010",
62 => "011010111Y1111000001101001001000",
63 => "11Y01101010010010110001010000010",
64 => "111001100110110110101000Y1010001",
65 => "011001101010101110101011Y1001111",
66 => "00010000000111101Y00110101101110",
67 => "10Y01110111111110101001011111111",
68 => "11000100011011001011Y11000111100",
69 => "00010000100001100000Y01000011011",
70 => "10000000101110101101100Y01010000",
71 => "11001010010011101010000Y11101011",
72 => "0010010010100100100001110000Y111",
73 => "101101101110001100000001000Y0011",
74 => "1001101100000110011101101011Y000",
75 => "110111Y0000000010111111111001111",
76 => "100100001Y1101010011100110000101",
77 => "11010000000101111Y11011010100101",
78 => "001100010101110000100101110Y1111",
79 => "100010101Y0010001000010111111100",
80 => "01Y01111010001001101100001001001",
81 => "0001011100000010111111011101111Y",
82 => "1001Y001110011100011111001000001",
83 => "100101101001000001Y0001001101001",
84 => "100101010101110000101011011011Y0",
85 => "1010110Y111110111111110001101110",
86 => "1111110110Y110101011000010101101",
87 => "101110101Y1011111011000000101111",
88 => "0100Y000111000011100101101010010",
89 => "1101010001010110101Y101111010001",
others => "00000000000000000000000000000000"),
(
0 => "0001111111100Y11000101Y100101001",
1 => "1100101Y0100010111000010000Y1000",
2 => "1100000010100111110YY10010101110",
3 => "1Y111Y10010010000101011011000010",
4 => "0110111011000110011100011001Y11Y",
5 => "001101Y111100101100001000111111Y",
6 => "0110Y00110010001100011000011100Y",
7 => "001100Y0110Y10011110110001000000",
8 => "110101Y111Y000111010000100100100",
9 => "000Y0101Y01111000001101110100011",
10 => "01101YY1110001101000110010000101",
11 => "10111111111010110000100Y1Y111011",
12 => "11011001Y001100111111001010Y1000",
13 => "0Y000011001100101111100Y11100111",
14 => "1010010111100111Y0000011Y0110011",
15 => "000Y0110111001Y11000101000111001",
16 => "001111010100111010101001Y0Y01011",
17 => "10011010101Y10010Y10010101111011",
18 => "10000000011011101Y1001101011Y011",
19 => "1111001110Y01Y110100010100001111",
20 => "111000011Y00111011010Y1001010110",
21 => "00Y011001011101000Y0001111010100",
22 => "100Y111Y101110100010011101100001",
23 => "001011100Y1001110010101Y01101001",
24 => "00011110110011101001YY0000101111",
25 => "110110000110000111101110Y110Y101",
26 => "110011000111100111111001100YY111",
27 => "1100110Y10011110110100000Y010100",
28 => "110110110000100101000Y1001001Y11",
29 => "110000010011011111001001Y011Y000",
30 => "01110100011011100101000Y0101110Y",
31 => "1101Y01001Y000101101111011100010",
32 => "110000100110010111110111100Y0010",
33 => "1100000011Y100101100001001110101",
34 => "1011110Y0000Y0110011101101111111",
35 => "01000011010010010010010Y0010011Y",
36 => "10000001111Y0001100010Y110111010",
37 => "10100001000000111Y11100001011Y01",
38 => "11101001110001100Y1110Y100110000",
39 => "00110001101111Y011Y0100000010111",
40 => "10000Y0001000Y010011100010000100",
41 => "0111111110110010Y0011001100110Y0",
42 => "1111001100010011011Y010Y10100000",
43 => "11111010Y0111111110Y101010101100",
44 => "110001101101100Y00000Y0101111110",
45 => "11100001110000Y010110001001000Y0",
46 => "111Y011000100011000010011001Y111",
47 => "1Y10100010001011110Y110110101111",
48 => "10011Y01110001Y11000001110100111",
49 => "01Y0011Y110110101100100010010100",
50 => "101101Y10111110011Y1101010100001",
51 => "001000000100011Y0Y00011100011110",
52 => "010110011110001100YY011001001100",
53 => "01110000000110001101000Y0000100Y",
54 => "1000000110011101Y101010100Y11111",
55 => "01001001101110011001Y11101001Y10",
56 => "10111011000001Y00100001000Y00000",
57 => "11001Y01111110101110000100Y01110",
58 => "111101Y1011010010001101Y00110100",
59 => "001000000101Y001110111010Y110010",
60 => "111100111Y0100Y11001010111100001",
61 => "101101100110Y01101010Y1101001100",
62 => "01001100111101101Y0110Y001100010",
63 => "000011101Y0000111101Y11001010111",
64 => "00001001010101000Y11Y11000101001",
65 => "0010010Y110001000Y01100101010101",
66 => "0100001011Y01011100110100Y101010",
67 => "000110101Y00101010Y1011000010100",
68 => "101100111111Y0101101Y00111011111",
69 => "10Y101110010000101101111000Y0100",
70 => "10001110001Y011001100Y0100110111",
71 => "00101Y1111110Y010100011000101101",
72 => "10111Y01Y00101010010101111000010",
73 => "011Y11Y0100101010000001010001001",
74 => "0Y1100101100011011101000100Y0011",
75 => "01000010110100010100110Y1100101Y",
76 => "11000010Y1011010000001100Y100010",
77 => "01Y00110101111101010000100Y00000",
78 => "000000000011100Y100101001010010Y",
79 => "011000Y1111000101001010Y10100001",
others => "00000000000000000000000000000000"),
(
0 => "010001100Y0010110111000001Y1Y100",
1 => "1111Y101110000011101001000Y00Y00",
2 => "011110Y1100111011110100100Y01010",
3 => "0Y111110110010001Y00011001010Y01",
4 => "1100Y01Y011Y01010011101001100011",
5 => "110Y01Y100011001Y000000010010001",
6 => "10Y10Y01Y10100101100001011010111",
7 => "100101000Y0001010Y111Y1001011010",
8 => "001011011001110100001010001YYY10",
9 => "1Y00010100010011Y1100110Y1110110",
10 => "1101001Y1100010011Y01100100110Y1",
11 => "0000Y11001001Y0011010Y1011111001",
12 => "101010011100010110Y11101Y1Y00110",
13 => "11000Y100100011Y0111100010010Y10",
14 => "111111100001100110YY101Y11000111",
15 => "1010010Y001101YY1111111100011111",
16 => "10000Y1110110Y10110110010100111Y",
17 => "1110000Y00Y1110100101111101Y1101",
18 => "01000011Y100001000Y1Y10101100011",
19 => "0Y111000111000101Y110111100Y1010",
20 => "010100011010101001001101Y00Y101Y",
21 => "00010100Y10100111Y00010001110011",
22 => "01110010100101011Y00Y110111Y0110",
23 => "00Y10000110101001011100Y01110001",
24 => "1010Y00Y00011Y000111011001111001",
25 => "0Y0101Y11000111100001100Y0000111",
26 => "100011Y1111001Y100Y0110000011110",
27 => "010Y1111101011100011101Y1110101Y",
28 => "001011000111111011000Y100Y0010Y1",
29 => "1011111011001011110110Y0011Y1011",
30 => "111101001Y10011111100010Y1010Y01",
31 => "100Y11Y1000001111000Y10100001011",
32 => "1111Y1101000110000010000Y11001Y0",
33 => "1100111011Y00100101Y10101010Y000",
34 => "111010110100100101Y010Y010011Y10",
35 => "011001100001101010Y10011Y1Y00111",
36 => "101100Y10101010000010001Y011001Y",
37 => "0011100101YY1010011110010000001Y",
38 => "10101110Y0101011Y10000Y110100110",
39 => "0110011Y110Y10111Y01000010110000",
40 => "0000010010100000111Y01Y0011101Y1",
41 => "0110011111Y11111Y000101010100110",
42 => "10001101110101Y01Y01000010Y01111",
43 => "0010001110Y01101000010101100Y001",
44 => "01Y01010Y1101Y001101111101111010",
45 => "101011001101011Y001111010001100Y",
46 => "1110Y1111Y1110101001001100011011",
47 => "111000100001Y011010010111Y001Y10",
48 => "1101010101111010000110Y1001Y101Y",
49 => "01Y0000Y10100Y100101111100101011",
50 => "101011111Y1100011Y0010Y000100100",
51 => "10100101111110110Y101010Y110001Y",
52 => "11111010YYY110000001000101000100",
53 => "01100Y0011Y1010101Y0110101101001",
54 => "101100111100001010Y101000YY01000",
55 => "0Y101010011011100101000110Y1010Y",
56 => "001110011101001001Y101Y01Y000111",
57 => "11010111110Y010111010101Y111Y010",
58 => "00Y00110100001110110010000101Y1Y",
59 => "100Y00101001Y111111101111101111Y",
60 => "110YY0100100000010001110011Y1010",
61 => "10100010Y011000Y10100Y1010011100",
62 => "100101100Y011100001110110Y11Y011",
63 => "0YY110100101111111110Y1011111101",
64 => "101Y111001111011000011010011YY00",
65 => "0101Y0110Y11111101Y0010001010000",
66 => "001101100000110Y000101Y1000100Y0",
67 => "01101Y1Y0100100111100000000Y0001",
68 => "1011100111001Y01011111011Y111001",
69 => "1Y01010000111111100000101110Y1Y0",
others => "00000000000000000000000000000000"),
(
0 => "1011111Y0Y1011001101Y11000001010",
1 => "10Y1010111Y1101111001Y1Y00010010",
2 => "111100Y1110110100Y00011110Y10111",
3 => "10Y01001101011Y11Y101001011Y0100",
4 => "10100Y10Y0011010001110Y11101Y000",
5 => "11Y0Y01001101000101100010000Y00Y",
6 => "1001100110Y01011Y010110Y1011Y110",
7 => "1010Y10101000Y1111001Y1001100Y10",
8 => "0110000101011YY100111000Y101Y110",
9 => "100Y00110100101011011Y110Y10111Y",
10 => "1000000011100YY0Y01110110Y000111",
11 => "100Y11001Y0000000110101101Y001Y1",
12 => "1Y101Y111000001Y1010111101111010",
13 => "00000111101Y00000100000Y11001Y11",
14 => "010101YY10101Y0Y0011010001100010",
15 => "10111101001Y101101000Y00011Y00Y0",
16 => "11101010Y110111001000101Y1Y11Y10",
17 => "1Y10Y0000110YY001001011101000011",
18 => "0Y01Y0Y0110010000001Y01001100000",
19 => "10Y0011010000110111YY001Y0000110",
20 => "1010110YY000010100101110101Y0Y01",
21 => "11000000011001Y1101Y0Y100011101Y",
22 => "1000110Y110110010Y100111110Y11Y0",
23 => "1111Y00Y10011101110110111Y11Y000",
24 => "00Y11011100010011Y1Y1110010100Y1",
25 => "0101100111001101Y1110Y0011110YY1",
26 => "1100001110110011Y0111Y110010Y00Y",
27 => "1Y1Y111Y010Y10101100111011010101",
28 => "10001011Y1010011101Y11Y101100Y01",
29 => "1Y0010110000011100Y0Y00Y00001111",
30 => "00000Y1101100Y11Y0101001001101Y1",
31 => "101000010100100Y0Y010000001101YY",
32 => "010001Y1011010001111011010Y11Y0Y",
33 => "01011011100011Y0Y101111Y11100111",
34 => "1Y1Y1Y101011Y1111000101111101111",
35 => "0Y01101Y11YY10010000010011010110",
36 => "110001Y010YY10101Y01110110100100",
37 => "101000110Y100Y00Y0Y0000001000010",
38 => "10010Y01Y11000110100010101011YY1",
39 => "11101110Y01101Y01110101Y01011101",
40 => "0Y110010Y01100Y1011101Y101001010",
41 => "01001010101Y1Y101111Y10101101001",
42 => "10110Y100Y100Y11011000101110111Y",
43 => "01Y1101101010Y1110100011110011Y1",
44 => "10010110111001001100100010YY10Y1",
45 => "1110010011001Y10Y10Y1Y0000100111",
46 => "0111Y0000100YY1110010001001Y0000",
47 => "01Y1010011111001010011011Y1Y0Y01",
48 => "101110101YY01001Y00000111100Y000",
49 => "100011Y10Y1Y100000000111001101Y1",
50 => "0101Y11100101000Y010010111Y1000Y",
51 => "001001Y011111Y0110110100011Y01Y1",
52 => "010111111000001100001010001Y0Y11",
53 => "0110Y001011Y101001011000010Y10Y1",
54 => "010010101101YY11100101001111Y0Y1",
55 => "00Y1111101Y010111111011Y01Y01110",
56 => "110000110011YY101Y101000010Y0110",
57 => "00000001YY011100001Y11111110Y000",
58 => "11001011111Y0111Y100Y1100100Y111",
59 => "101110101101111Y00Y0001110000Y0Y",
others => "00000000000000000000000000000000"),
(
0 => "0001Y01101111011Y100Y0000010YY10",
1 => "1011Y0Y0110101011Y1101010Y100100",
2 => "1Y0010010111Y10101000Y110Y11Y001",
3 => "1011100Y0101111Y101011Y001Y0101Y",
4 => "0001011YY0000111Y01011111111Y101",
5 => "01Y0YY11011001101000110YY1100101",
6 => "01Y0100010101Y1100Y1100000Y0110Y",
7 => "10Y010000011101YY0010100001YY010",
8 => "000Y00Y0011Y11000001Y10011010Y01",
9 => "011Y00100Y1111100100001YY000011Y",
10 => "1YY0010111Y11Y110Y00110101000011",
11 => "100000YY0110001110YY11100101Y010",
12 => "11001010111011010YY1010100YY11Y0",
13 => "10Y110Y1101111001000111000Y10100",
14 => "00Y110111010Y0Y01110001YY0001100",
15 => "1010000101110Y111110010Y0YY10011",
16 => "010110000100101Y1Y0110Y110Y001Y1",
17 => "0001000001000Y100111011Y00YY00Y1",
18 => "101Y101100111Y111100Y10Y10Y11111",
19 => "11Y1101110101101010YY001001Y1Y11",
20 => "011101Y110110010Y10Y00010111Y01Y",
21 => "1100001YY001Y000Y0000110011Y1111",
22 => "100Y0Y0010001Y001Y1110Y000010100",
23 => "11001011Y0000Y00Y1100000011Y1101",
24 => "010Y01111Y0111YY000000001Y010100",
25 => "1Y01110000000100Y10Y010Y11000Y11",
26 => "01010Y00001110YYYY00111011111010",
27 => "000Y110Y0111110100001Y11Y0110000",
28 => "11Y1111100Y011110100Y10110Y0Y111",
29 => "00011110YY1Y1000011011100001Y01Y",
30 => "1Y00010Y101Y11010111Y1000Y100010",
31 => "101Y000110101000Y0Y0Y1101Y100110",
32 => "1001110Y00Y1Y0Y110010100011001Y1",
33 => "111011011Y0011100YY0001Y10Y01111",
34 => "1000101Y0Y01011YY00Y011111000110",
35 => "1000000111Y0Y010010Y10101000Y001",
36 => "00Y1101010000Y11000111Y00Y010011",
37 => "00010011111100Y11011110YY0111Y00",
38 => "0Y001010000Y0011Y01001000001YY10",
39 => "0Y11Y00001111101101000YY1Y001000",
40 => "101Y10111YY101010001Y0110Y110101",
41 => "001Y001001001111Y1Y0001Y01010011",
42 => "01111YY0Y110000010100001Y0011100",
43 => "100110001001Y10000111010Y0111YYY",
44 => "1000000000110Y011Y001110Y01Y0010",
45 => "0101011Y111010111110Y1YY1111110Y",
46 => "1001Y110110101YY111001010100Y110",
47 => "000101001011011111Y1Y001101111YY",
48 => "11110110Y1Y0110YY1Y0001101101010",
49 => "0Y0Y10111111Y0100001Y11100000Y00",
others => "00000000000000000000000000000000"),
(
0 => "1Y11110011001Y00Y011101Y11110Y01",
1 => "11Y010000Y110Y10Y010111010100Y1Y",
2 => "0011Y11Y011Y10110011101010Y0YY11",
3 => "00Y1Y1Y1Y1110011YY11011100000011",
4 => "11000111Y11Y11111Y0Y10000101YY01",
5 => "1010110011Y1010Y10Y0101Y001Y101Y",
6 => "0010110001Y010Y111Y010100Y1Y101Y",
7 => "1111Y10Y01111Y111010Y0Y10011Y010",
8 => "1000000Y100011Y1001100010Y0Y10YY",
9 => "00011Y01101Y10Y0111101Y00111110Y",
10 => "11Y0Y101001010Y10111Y1111101YY00",
11 => "1Y11110Y00Y101011Y10101000101Y0Y",
12 => "1Y0111Y11000Y0Y0Y101001Y00001100",
13 => "0100101Y111Y1100110101Y00Y10Y000",
14 => "01101110Y1000YY001001Y000Y000000",
15 => "01Y1101Y001000Y101Y1Y1Y111101001",
16 => "00Y100000Y1110100011Y1Y1Y110Y101",
17 => "01Y00Y1Y111000Y0011001111Y1Y1010",
18 => "11011100010010Y001Y0001YY00Y0100",
19 => "010YYY1001111001110YY100Y0101111",
20 => "010Y10Y0Y000000110Y01001011Y1101",
21 => "01110110111Y000010001YYY0Y011010",
22 => "00Y010001Y01110Y10Y1Y010101Y1001",
23 => "1Y0011000101Y0100Y111Y1110010001",
24 => "011111111Y0010Y01YY110Y1110000Y1",
25 => "110Y111110000Y01110100Y000Y110Y1",
26 => "0101110011111Y01YY110Y1000110YY0",
27 => "010Y0YYY1Y011100111010000010Y001",
28 => "011101Y01Y01Y010010Y100011Y111Y1",
29 => "01110100111Y0Y000111001Y10YY1000",
30 => "11Y10000101001000Y101110YYY10111",
31 => "11Y0010Y11Y1Y0010111111001Y0Y101",
32 => "1Y101100001Y11111101Y001Y1010Y10",
33 => "10Y111Y11Y0Y0111111011100Y00Y011",
34 => "100000Y001Y00100Y10010Y1YY001111",
35 => "01YY0Y111Y000001000000Y101110Y10",
36 => "01001001100101Y1Y00100Y0Y0011Y1Y",
37 => "0Y000101011YY01111000101Y00Y0000",
38 => "101Y0100Y010111010Y1Y1010Y1100Y0",
39 => "01Y0Y0100100110Y00010000Y1010101",
others => "00000000000000000000000000000000"),
(
0 => "0Y1Y0001Y01011011110001010Y00Y1Y",
1 => "10001YYY00101010Y01011100010Y0YY",
2 => "0Y01111Y010Y1Y10000110000Y11Y001",
3 => "1101Y00Y01Y101Y10Y0000001001Y101",
4 => "110101Y111100110Y1000Y0Y110Y000Y",
5 => "0Y00101111101000Y11YY000Y0011100",
6 => "0010Y1110Y101100111101101Y1001YY",
7 => "001101101001YY110Y0YY10100Y10100",
8 => "1Y0111Y0111Y010Y11000Y1Y0Y110010",
9 => "11YY11000Y110YY0100Y0110Y0100111",
10 => "001100Y111YYY01100Y110Y1011000Y1",
11 => "1Y1Y01010011Y1111Y01Y11101Y0101Y",
12 => "0001Y1011Y010000100000Y0Y0101YY0",
13 => "1001100001101YY100YY101001Y01Y0Y",
14 => "10011100YY10001Y1Y1Y1Y101000110Y",
15 => "1110110Y0111011YY0Y10Y001Y111011",
16 => "0Y100Y010011100Y00YY0101001Y100Y",
17 => "00010YY01YY111010Y0010Y000Y11100",
18 => "11Y0Y1Y1Y111010011011111001YY11Y",
19 => "0YY101Y110000000100Y111Y01Y111Y1",
20 => "0001YY01100110Y00Y00Y1011111100Y",
21 => "0101Y00YY01010Y111Y11Y1011010110",
22 => "11Y0000100111111010Y01Y10001YYY0",
23 => "00111YY10Y110100000Y00Y1Y100111Y",
24 => "01001100Y0YY1111Y0111Y01Y1101001",
25 => "111010110Y1Y11YY001Y1110000Y1Y11",
26 => "01000Y010110100YY1010Y0001Y01Y0Y",
27 => "1Y01Y01011111000110Y1Y00Y01111Y1",
28 => "010Y111011Y0YY01Y01001111YY11100",
29 => "10Y0000Y10011Y0010Y1011Y1YY00111",
others => "00000000000000000000000000000000"),
(
0 => "01001YY010Y11101110010Y10Y1YY1Y0",
1 => "1000YY0Y001Y1Y111001Y0000001Y001",
2 => "0Y0Y1YY110Y0Y100Y101011101001000",
3 => "1Y1101Y1111Y11001111Y001100YYYY0",
4 => "1010Y111Y1100Y0100100010Y001YY1Y",
5 => "0001000Y111YY1000101YYY01101011Y",
6 => "1101Y101010011000Y1Y01Y00Y1110YY",
7 => "0Y01Y110100Y010YY001110Y001101Y0",
8 => "1Y11Y1110Y0Y110001YYY0100111Y001",
9 => "10011Y11Y10Y0YY001Y1110011100Y10",
10 => "10Y0101Y10Y0111001111YY00110Y000",
11 => "011YY01111YY01Y01Y1101000110Y011",
12 => "1Y10110Y1100Y1001Y1Y11Y1101YY010",
13 => "0Y1Y1011YY0101000000110YY01YY100",
14 => "0Y1YY1011111Y11110Y11Y0YY0001110",
15 => "00001Y00111Y00001011Y1011YY0Y010",
16 => "001YY010011Y0Y010011101111Y1Y010",
17 => "111Y000001Y0Y110001Y0010011Y0Y00",
18 => "1111110YY0Y010100Y111Y110Y01Y011",
19 => "01111Y10Y1001Y111011Y011Y0Y0Y1Y1",
others => "00000000000000000000000000000000"),
(
0 => "10Y0100100Y1Y0YY11Y1Y00Y11000Y11",
1 => "010YYY00Y1Y010Y100000011Y111011Y",
2 => "0Y01111Y10101Y010YY0100Y01YY0011",
3 => "001YY0001Y0110Y1111010Y00011Y001",
4 => "00010YY0YY10Y00YY001Y101Y1001011",
5 => "10Y0Y110Y1000000Y1101Y10YY11Y010",
6 => "0Y000Y1Y00Y01Y101100Y0Y01001111Y",
7 => "0001101Y0Y100YYY0001100001Y1110Y",
8 => "1Y101Y1110Y0101110Y10Y0Y0Y0YY110",
9 => "01011YY011Y110YYY111YY1000001010",
others => "00000000000000000000000000000000")
);
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;