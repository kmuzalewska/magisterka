library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
library xil_defaultlib;
use xil_defaultlib.types.all;

package data_to_tcam is

constant DATA_TO_TCAM_CONST : TCAM_ARRAY_3D :=
(
(
0 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
1 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
2 => ("00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
3 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01"),
4 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
5 => ("01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01"),
6 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
7 => ("01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00"),
8 => ("01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
9 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00"),
10 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
11 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01"),
12 => ("00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
13 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00"),
14 => ("01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01"),
15 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
16 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01"),
17 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
18 => ("01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
19 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
20 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
21 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00"),
22 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
23 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
24 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
25 => ("00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01"),
26 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00"),
27 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
28 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
29 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00"),
30 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
31 => ("01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00"),
32 => ("00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
33 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
34 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
35 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00"),
36 => ("00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
37 => ("00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
38 => ("01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
39 => ("01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
40 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01"),
41 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00"),
42 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
43 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
44 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
45 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
46 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00"),
47 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01"),
48 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
49 => ("00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01"),
50 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
51 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
52 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
53 => ("01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
54 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01"),
55 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
56 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
57 => ("00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00"),
58 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
59 => ("01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01"),
60 => ("01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01"),
61 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01"),
62 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
63 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
64 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
65 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
66 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
67 => ("00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
68 => ("01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
69 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00"),
70 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01"),
71 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01"),
72 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01"),
73 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
74 => ("00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01"),
75 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
76 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01"),
77 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01"),
78 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01"),
79 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00"),
80 => ("00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
81 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
82 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
83 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00"),
84 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01"),
85 => ("00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
86 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
87 => ("00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00"),
88 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
89 => ("01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00"),
90 => ("00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00"),
91 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00"),
92 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00"),
93 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00"),
94 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
95 => ("00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
96 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
97 => ("00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01"),
98 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01"),
99 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01"),
100 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01"),
101 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
102 => ("00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01"),
103 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
104 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01"),
105 => ("01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
106 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
107 => ("01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
108 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01"),
109 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
110 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
111 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01"),
112 => ("00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01"),
113 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00"),
114 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
115 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01"),
116 => ("01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
117 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00"),
118 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
119 => ("01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
120 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01"),
121 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01"),
122 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00"),
123 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
124 => ("01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
125 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00"),
126 => ("00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
127 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
128 => ("01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
129 => ("00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00"),
130 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01"),
131 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
132 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01"),
133 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
134 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
135 => ("01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01"),
136 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
137 => ("01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00"),
138 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
139 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01"),
140 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01"),
141 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
142 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
143 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01"),
144 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
145 => ("00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01"),
146 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00"),
147 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
148 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
149 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
150 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01"),
151 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
152 => ("01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
153 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01"),
154 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00"),
155 => ("01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00"),
156 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01"),
157 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01"),
158 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
159 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
160 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
161 => ("01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
162 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
163 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
164 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00"),
165 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01"),
166 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
167 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01"),
168 => ("00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01"),
169 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01"),
170 => ("00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
171 => ("01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01"),
172 => ("01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01"),
173 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01"),
174 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00"),
175 => ("00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
176 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
177 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
178 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01"),
179 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
180 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
181 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
182 => ("00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
183 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
184 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
185 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
186 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
187 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
188 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
189 => ("01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
190 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
191 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
192 => ("00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
193 => ("00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01"),
194 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
195 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
196 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
197 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
198 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
199 => ("00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
200 => ("01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00"),
201 => ("01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01"),
202 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01"),
203 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00"),
204 => ("01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
205 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00"),
206 => ("01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00"),
207 => ("01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
208 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
209 => ("01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00"),
210 => ("00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
211 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00"),
212 => ("01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00"),
213 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01"),
214 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
215 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
216 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
217 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
218 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00"),
219 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
220 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00"),
221 => ("00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
222 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00"),
223 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
224 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
225 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00"),
226 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
227 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01"),
228 => ("01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
229 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00"),
230 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00"),
231 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
232 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
233 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01"),
234 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
235 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
236 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
237 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
238 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
239 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
240 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
241 => ("00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01"),
242 => ("01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00"),
243 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00"),
244 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00"),
245 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01"),
246 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01"),
247 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
248 => ("01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
249 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
250 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
251 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
252 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
253 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
254 => ("01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01"),
255 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00"),
256 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
257 => ("01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00"),
258 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00"),
259 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01"),
260 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00"),
261 => ("01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01"),
262 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
263 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01"),
264 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
265 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01"),
266 => ("01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
267 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
268 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
269 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
270 => ("00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00"),
271 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
272 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
273 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
274 => ("01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
275 => ("01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00"),
276 => ("01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01"),
277 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00"),
278 => ("00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01"),
279 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
280 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
281 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
282 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
283 => ("01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
284 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
285 => ("01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
286 => ("00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
287 => ("01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
288 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
289 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01"),
290 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
291 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
292 => ("01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
293 => ("01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
294 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
295 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
296 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
297 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00"),
298 => ("00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
299 => ("01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
300 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01"),
301 => ("01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01"),
302 => ("01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01"),
303 => ("00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
304 => ("00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
305 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
306 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00"),
307 => ("00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00"),
308 => ("01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
309 => ("01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00"),
310 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
311 => ("00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00"),
312 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
313 => ("01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01"),
314 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
315 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
316 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
317 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
318 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01"),
319 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01"),
320 => ("01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
321 => ("00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01"),
322 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01"),
323 => ("00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
324 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
325 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
326 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
327 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
328 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
329 => ("00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
330 => ("01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
331 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
332 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
333 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01"),
334 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
335 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01"),
336 => ("01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
337 => ("01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01"),
338 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
339 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
340 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
341 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
342 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
343 => ("01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00"),
344 => ("01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01"),
345 => ("01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01"),
346 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
347 => ("00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01"),
348 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00"),
349 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
350 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00"),
351 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
352 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
353 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
354 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
355 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
356 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
357 => ("00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00"),
358 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
359 => ("01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00"),
360 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
361 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
362 => ("01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01"),
363 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01"),
364 => ("01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
365 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
366 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
367 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01"),
368 => ("01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
369 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
370 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01"),
371 => ("00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01"),
372 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01"),
373 => ("01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00"),
374 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01"),
375 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
376 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00"),
377 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01"),
378 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01"),
379 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
380 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
381 => ("01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
382 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
383 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00"),
384 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
385 => ("00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01"),
386 => ("01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
387 => ("00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00"),
388 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
389 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00"),
390 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01"),
391 => ("01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
392 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
393 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
394 => ("01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00"),
395 => ("00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00"),
396 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
397 => ("01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
398 => ("01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01"),
399 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00"),
400 => ("00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
401 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01"),
402 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
403 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
404 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00"),
405 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
406 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01"),
407 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
408 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
409 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
410 => ("01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
411 => ("01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01"),
412 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
413 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
414 => ("01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
415 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
416 => ("01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01"),
417 => ("01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00"),
418 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
419 => ("00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
420 => ("01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00"),
421 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00"),
422 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
423 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01"),
424 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
425 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
426 => ("01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00"),
427 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00"),
428 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
429 => ("01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
430 => ("00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
431 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01"),
432 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00"),
433 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00"),
434 => ("01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01"),
435 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
436 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
437 => ("01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
438 => ("00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01"),
439 => ("00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
440 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00"),
441 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
442 => ("01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
443 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
444 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
445 => ("01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
446 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
447 => ("01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00"),
448 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01"),
449 => ("01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01"),
450 => ("00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
451 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00"),
452 => ("01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00"),
453 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
454 => ("01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
455 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00"),
456 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01"),
457 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01"),
458 => ("00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
459 => ("00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
460 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00"),
461 => ("01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
462 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
463 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
464 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
465 => ("00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
466 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
467 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
468 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
469 => ("01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
470 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
471 => ("01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00"),
472 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01"),
473 => ("00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
474 => ("00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
475 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01"),
476 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
477 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
478 => ("00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01"),
479 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
480 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"),
481 => ("00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
482 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01"),
483 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
484 => ("01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
485 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
486 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01"),
487 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00"),
488 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
489 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
490 => ("00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01"),
491 => ("01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
492 => ("00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
493 => ("01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
494 => ("01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00"),
495 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01"),
496 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
497 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01"),
498 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
499 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01")),
(
0 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00"),
1 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01"),
2 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01"),
3 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01"),
4 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11"),
5 => ("00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
6 => ("00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00"),
7 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01"),
8 => ("01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01"),
9 => ("00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00"),
10 => ("01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
11 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
12 => ("00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01"),
13 => ("00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "00"),
14 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01"),
15 => ("01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01"),
16 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01"),
17 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
18 => ("00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00"),
19 => ("01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
20 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01"),
21 => ("00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
22 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00"),
23 => ("01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
24 => ("00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
25 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
26 => ("01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01"),
27 => ("01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01"),
28 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
29 => ("01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
30 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00"),
31 => ("00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00"),
32 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
33 => ("01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00"),
34 => ("00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
35 => ("01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11"),
36 => ("00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00"),
37 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01"),
38 => ("01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
39 => ("01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00"),
40 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
41 => ("01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01"),
42 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00"),
43 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00"),
44 => ("00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00"),
45 => ("01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01"),
46 => ("00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
47 => ("00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
48 => ("00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
49 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01"),
50 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
51 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00"),
52 => ("00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00"),
53 => ("00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00"),
54 => ("00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
55 => ("01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
56 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01"),
57 => ("01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01"),
58 => ("00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01"),
59 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01"),
60 => ("01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "00"),
61 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01"),
62 => ("00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
63 => ("01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00"),
64 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00"),
65 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01"),
66 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00"),
67 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
68 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
69 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01"),
70 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
71 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01"),
72 => ("00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01"),
73 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01"),
74 => ("01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
75 => ("00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
76 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
77 => ("01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
78 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
79 => ("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00"),
80 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01"),
81 => ("01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
82 => ("01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
83 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
84 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
85 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00"),
86 => ("00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01"),
87 => ("01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
88 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01"),
89 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01"),
90 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01"),
91 => ("01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
92 => ("01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00"),
93 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01"),
94 => ("00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01"),
95 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
96 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00"),
97 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
98 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00"),
99 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
100 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
101 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01"),
102 => ("00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
103 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00"),
104 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
105 => ("01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
106 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
107 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01"),
108 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
109 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
110 => ("01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
111 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01"),
112 => ("01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01"),
113 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01"),
114 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01"),
115 => ("01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
116 => ("01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01"),
117 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
118 => ("01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
119 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00"),
120 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01"),
121 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00"),
122 => ("01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11"),
123 => ("01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
124 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01"),
125 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00"),
126 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
127 => ("01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01"),
128 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
129 => ("00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01"),
130 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00"),
131 => ("01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
132 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11"),
133 => ("00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
134 => ("00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00"),
135 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01"),
136 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
137 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
138 => ("01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00"),
139 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01"),
140 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01"),
141 => ("00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
142 => ("01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
143 => ("01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
144 => ("01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
145 => ("00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01"),
146 => ("00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01"),
147 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01"),
148 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
149 => ("00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00"),
150 => ("00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00"),
151 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00"),
152 => ("01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
153 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01"),
154 => ("01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
155 => ("00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01"),
156 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00"),
157 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00"),
158 => ("00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
159 => ("01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
160 => ("01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00"),
161 => ("00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
162 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00"),
163 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01"),
164 => ("00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01"),
165 => ("01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
166 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
167 => ("01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
168 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11"),
169 => ("00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
170 => ("00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11"),
171 => ("00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
172 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
173 => ("00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
174 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
175 => ("01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
176 => ("00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
177 => ("00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00"),
178 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00"),
179 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00"),
180 => ("01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01"),
181 => ("00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00"),
182 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00"),
183 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00"),
184 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00"),
185 => ("00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00"),
186 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
187 => ("00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00"),
188 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00"),
189 => ("01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01"),
190 => ("01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00"),
191 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00"),
192 => ("01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
193 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
194 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01"),
195 => ("00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01"),
196 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01"),
197 => ("01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
198 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01"),
199 => ("01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
200 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01"),
201 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01"),
202 => ("00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
203 => ("01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00"),
204 => ("00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
205 => ("01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
206 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00"),
207 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01"),
208 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01"),
209 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
210 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01"),
211 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
212 => ("00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01"),
213 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01"),
214 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00"),
215 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
216 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
217 => ("01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
218 => ("00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00"),
219 => ("00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00"),
220 => ("01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
221 => ("00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01"),
222 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00"),
223 => ("01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00"),
224 => ("01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01"),
225 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00"),
226 => ("01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00"),
227 => ("00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00"),
228 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
229 => ("01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01"),
230 => ("00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
231 => ("00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01"),
232 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01"),
233 => ("01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00"),
234 => ("00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00"),
235 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01"),
236 => ("01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
237 => ("01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
238 => ("01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01"),
239 => ("01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00"),
240 => ("00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
241 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
242 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00"),
243 => ("00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
244 => ("00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00"),
245 => ("00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
246 => ("01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00"),
247 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01"),
248 => ("01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
249 => ("01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01"),
250 => ("00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
251 => ("01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01"),
252 => ("01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
253 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
254 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01"),
255 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01"),
256 => ("01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
257 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01"),
258 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "01"),
259 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
260 => ("01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01"),
261 => ("00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
262 => ("00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00"),
263 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01"),
264 => ("00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
265 => ("01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
266 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00"),
267 => ("00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
268 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00"),
269 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
270 => ("00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
271 => ("01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00"),
272 => ("01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "00"),
273 => ("00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00"),
274 => ("00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
275 => ("01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01"),
276 => ("01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01"),
277 => ("00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00"),
278 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
279 => ("01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00"),
280 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
281 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
282 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
283 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
284 => ("00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00"),
285 => ("01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
286 => ("01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00"),
287 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00"),
288 => ("00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
289 => ("00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
290 => ("01", "00", "11", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01"),
291 => ("00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01"),
292 => ("01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01"),
293 => ("01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
294 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00"),
295 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
296 => ("01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
297 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00"),
298 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
299 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01"),
300 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00"),
301 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
302 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
303 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01"),
304 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
305 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
306 => ("00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01"),
307 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00"),
308 => ("01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
309 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11"),
310 => ("01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00"),
311 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
312 => ("00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
313 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00"),
314 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01"),
315 => ("01", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00"),
316 => ("01", "11", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
317 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
318 => ("00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
319 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
320 => ("01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01"),
321 => ("01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00"),
322 => ("00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
323 => ("01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01"),
324 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
325 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
326 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01"),
327 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00"),
328 => ("00", "00", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00"),
329 => ("00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00"),
330 => ("01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
331 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00"),
332 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00"),
333 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00"),
334 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00"),
335 => ("00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00"),
336 => ("00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00"),
337 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01"),
338 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00"),
339 => ("01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01"),
340 => ("00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
341 => ("01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01"),
342 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00"),
343 => ("01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01"),
344 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00"),
345 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00"),
346 => ("01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
347 => ("01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01"),
348 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01"),
349 => ("00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
350 => ("00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
351 => ("01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
352 => ("00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
353 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
354 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "00"),
355 => ("00", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01"),
356 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00"),
357 => ("01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
358 => ("00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
359 => ("01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01"),
360 => ("00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01"),
361 => ("01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00"),
362 => ("00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00"),
363 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00"),
364 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
365 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01"),
366 => ("01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
367 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00"),
368 => ("01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01"),
369 => ("01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00"),
370 => ("01", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00"),
371 => ("00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00"),
372 => ("01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
373 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01"),
374 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01"),
375 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00"),
376 => ("01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01"),
377 => ("00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
378 => ("00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01"),
379 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00"),
380 => ("00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
381 => ("01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
382 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00"),
383 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
384 => ("01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
385 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00"),
386 => ("00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01"),
387 => ("01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
388 => ("01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01"),
389 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
390 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00"),
391 => ("01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00"),
392 => ("00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
393 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00"),
394 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00"),
395 => ("00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00"),
396 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01"),
397 => ("01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
398 => ("00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01"),
399 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00"),
400 => ("01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
401 => ("00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
402 => ("00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00"),
403 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
404 => ("01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "00"),
405 => ("00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
406 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
407 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
408 => ("00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01"),
409 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
410 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00"),
411 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
412 => ("01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
413 => ("00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01"),
414 => ("01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00"),
415 => ("00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01"),
416 => ("00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
417 => ("01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
418 => ("00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01"),
419 => ("00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00"),
420 => ("00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
421 => ("01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
422 => ("00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
423 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
424 => ("00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00"),
425 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01"),
426 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01"),
427 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01"),
428 => ("01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
429 => ("00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
430 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00"),
431 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00"),
432 => ("01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
433 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01"),
434 => ("00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
435 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
436 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
437 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
438 => ("00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00"),
439 => ("01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
440 => ("01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00"),
441 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01"),
442 => ("01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01"),
443 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01"),
444 => ("01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01"),
445 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00"),
446 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
447 => ("00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01"),
448 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00"),
449 => ("00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00"),
450 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
451 => ("01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
452 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01"),
453 => ("00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01"),
454 => ("00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
455 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00"),
456 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00"),
457 => ("00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
458 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
459 => ("01", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00"),
460 => ("00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01"),
461 => ("01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
462 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00"),
463 => ("01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
464 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01"),
465 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
466 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01"),
467 => ("00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
468 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
469 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
470 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01"),
471 => ("00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
472 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
473 => ("01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00"),
474 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00"),
475 => ("01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
476 => ("00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
477 => ("00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
478 => ("01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01"),
479 => ("01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01"),
480 => ("01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01"),
481 => ("00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01"),
482 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00"),
483 => ("00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01"),
484 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00"),
485 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01"),
486 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
487 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00"),
488 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01"),
489 => ("01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11"),
490 => ("01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01"),
491 => ("01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00"),
492 => ("01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00"),
493 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00"),
494 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00"),
495 => ("01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
496 => ("01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00"),
497 => ("00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01"),
498 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
499 => ("01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00")),
(
0 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01"),
1 => ("00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01"),
2 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "01", "00"),
3 => ("01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
4 => ("00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01"),
5 => ("01", "00", "00", "00", "01", "00", "11", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
6 => ("00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
7 => ("01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01"),
8 => ("01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
9 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "11"),
10 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00"),
11 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00"),
12 => ("01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00", "00", "00"),
13 => ("01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
14 => ("00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01"),
15 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01"),
16 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01"),
17 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01"),
18 => ("00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
19 => ("00", "00", "00", "00", "11", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
20 => ("00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01"),
21 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01"),
22 => ("01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11"),
23 => ("01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
24 => ("01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11"),
25 => ("01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
26 => ("01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01"),
27 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "11", "00", "01", "01", "00"),
28 => ("01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01"),
29 => ("01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11"),
30 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
31 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00"),
32 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11"),
33 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "11", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01"),
34 => ("00", "01", "11", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
35 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
36 => ("00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11"),
37 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "11", "00"),
38 => ("01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "11", "01", "01", "01"),
39 => ("01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "11"),
40 => ("01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00"),
41 => ("00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01"),
42 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
43 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "00"),
44 => ("00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01"),
45 => ("01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01"),
46 => ("00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
47 => ("01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
48 => ("00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01"),
49 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
50 => ("00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11"),
51 => ("00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
52 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
53 => ("00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "11", "01", "00"),
54 => ("00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00"),
55 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01"),
56 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "11", "00", "01"),
57 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01"),
58 => ("01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
59 => ("00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
60 => ("00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01"),
61 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01"),
62 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01"),
63 => ("00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00"),
64 => ("00", "11", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
65 => ("01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11"),
66 => ("01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11"),
67 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00"),
68 => ("00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00"),
69 => ("01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01"),
70 => ("00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
71 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00"),
72 => ("01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
73 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01"),
74 => ("01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00"),
75 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00"),
76 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
77 => ("01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11"),
78 => ("00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
79 => ("00", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01"),
80 => ("01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01"),
81 => ("00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01"),
82 => ("01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01"),
83 => ("00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
84 => ("01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01"),
85 => ("01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00"),
86 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01"),
87 => ("00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01"),
88 => ("01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
89 => ("00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01"),
90 => ("00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
91 => ("01", "01", "01", "01", "00", "01", "11", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00"),
92 => ("00", "00", "01", "00", "11", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00"),
93 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
94 => ("01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01"),
95 => ("01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
96 => ("00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
97 => ("01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
98 => ("01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "11", "00", "01", "01"),
99 => ("01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
100 => ("00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
101 => ("01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
102 => ("00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01"),
103 => ("00", "01", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00"),
104 => ("01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "01"),
105 => ("01", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
106 => ("01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
107 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00"),
108 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00"),
109 => ("01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
110 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
111 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
112 => ("00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00"),
113 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00"),
114 => ("00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00"),
115 => ("01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
116 => ("00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01"),
117 => ("01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
118 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
119 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00"),
120 => ("01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01"),
121 => ("01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01"),
122 => ("00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00"),
123 => ("00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01"),
124 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "01", "01"),
125 => ("01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01"),
126 => ("01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00"),
127 => ("01", "01", "01", "11", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
128 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00"),
129 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00"),
130 => ("01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00"),
131 => ("00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00"),
132 => ("00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
133 => ("00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
134 => ("00", "00", "00", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01"),
135 => ("01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
136 => ("01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00"),
137 => ("01", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
138 => ("00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00"),
139 => ("00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "11"),
140 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
141 => ("00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
142 => ("00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01"),
143 => ("00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
144 => ("01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
145 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "00", "00"),
146 => ("01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00"),
147 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00"),
148 => ("00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
149 => ("00", "01", "00", "01", "00", "11", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
150 => ("00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00"),
151 => ("00", "00", "01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
152 => ("00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00"),
153 => ("01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00"),
154 => ("01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
155 => ("00", "11", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01"),
156 => ("01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01"),
157 => ("00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "01"),
158 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
159 => ("01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01"),
160 => ("01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00"),
161 => ("01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01"),
162 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11"),
163 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "11", "01", "01"),
164 => ("01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00"),
165 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
166 => ("00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00"),
167 => ("01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00"),
168 => ("00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01"),
169 => ("00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01"),
170 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00"),
171 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00"),
172 => ("00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01"),
173 => ("01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00"),
174 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00"),
175 => ("00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "11", "01", "01"),
176 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00"),
177 => ("00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00"),
178 => ("00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00"),
179 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "11", "01", "01", "01"),
180 => ("01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
181 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00"),
182 => ("00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11"),
183 => ("00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00"),
184 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00"),
185 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00"),
186 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00"),
187 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01"),
188 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00"),
189 => ("01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "01"),
190 => ("00", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00"),
191 => ("01", "01", "01", "11", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01"),
192 => ("00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01"),
193 => ("00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01"),
194 => ("00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00"),
195 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00"),
196 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00"),
197 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11"),
198 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11"),
199 => ("01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
200 => ("00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01"),
201 => ("00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00"),
202 => ("00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00"),
203 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00"),
204 => ("01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
205 => ("00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
206 => ("01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01"),
207 => ("00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01"),
208 => ("01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01"),
209 => ("00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01"),
210 => ("00", "00", "01", "01", "01", "11", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
211 => ("00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
212 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
213 => ("00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
214 => ("00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
215 => ("01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01"),
216 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01"),
217 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01"),
218 => ("01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00"),
219 => ("01", "01", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
220 => ("00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
221 => ("01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
222 => ("01", "00", "01", "00", "00", "01", "11", "00", "01", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
223 => ("00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01"),
224 => ("00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01"),
225 => ("01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01"),
226 => ("01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
227 => ("01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00"),
228 => ("00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11"),
229 => ("00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01"),
230 => ("00", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01"),
231 => ("00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
232 => ("01", "00", "11", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00"),
233 => ("01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11"),
234 => ("01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01"),
235 => ("00", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01"),
236 => ("01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00"),
237 => ("00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00"),
238 => ("00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01"),
239 => ("01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01"),
240 => ("01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
241 => ("00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00"),
242 => ("00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00"),
243 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00"),
244 => ("00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00"),
245 => ("01", "01", "01", "00", "00", "00", "01", "11", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00"),
246 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
247 => ("00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00"),
248 => ("00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01"),
249 => ("01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00"),
250 => ("00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
251 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00"),
252 => ("01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
253 => ("01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
254 => ("00", "01", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01"),
255 => ("01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01"),
256 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11"),
257 => ("00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01"),
258 => ("00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01"),
259 => ("00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00"),
260 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01"),
261 => ("01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00"),
262 => ("00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00"),
263 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01"),
264 => ("00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
265 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00"),
266 => ("00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00"),
267 => ("01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01"),
268 => ("01", "00", "00", "00", "00", "11", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01"),
269 => ("00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01"),
270 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
271 => ("01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
272 => ("00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00"),
273 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00"),
274 => ("00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
275 => ("00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
276 => ("01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11"),
277 => ("00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11"),
278 => ("01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00"),
279 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "11", "00"),
280 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "11", "00", "00", "00", "01", "00"),
281 => ("01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01"),
282 => ("01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
283 => ("01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
284 => ("00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
285 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
286 => ("00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00"),
287 => ("01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "11"),
288 => ("00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
289 => ("00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01"),
290 => ("00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
291 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01"),
292 => ("00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
293 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
294 => ("00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "01", "01"),
295 => ("00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01"),
296 => ("01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
297 => ("01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11"),
298 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "11", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
299 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01"),
300 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
301 => ("00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "00", "11", "00", "01"),
302 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11"),
303 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
304 => ("00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "11", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01"),
305 => ("00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01"),
306 => ("01", "01", "01", "01", "11", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01"),
307 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "11", "01", "00", "01"),
308 => ("01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00"),
309 => ("00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
310 => ("00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01"),
311 => ("01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01"),
312 => ("00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
313 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01"),
314 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11"),
315 => ("01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
316 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01"),
317 => ("01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00"),
318 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00"),
319 => ("00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00"),
320 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00"),
321 => ("01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01"),
322 => ("01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11"),
323 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "11", "00", "01", "01", "00", "01", "00", "00", "00"),
324 => ("01", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00"),
325 => ("01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
326 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01"),
327 => ("00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00"),
328 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
329 => ("01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00"),
330 => ("01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00"),
331 => ("00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01"),
332 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
333 => ("00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01"),
334 => ("00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01"),
335 => ("01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "00"),
336 => ("00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01"),
337 => ("01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01"),
338 => ("01", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00"),
339 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00"),
340 => ("00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01"),
341 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00"),
342 => ("01", "00", "01", "01", "11", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01"),
343 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00"),
344 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01"),
345 => ("01", "00", "00", "01", "00", "01", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01"),
346 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00"),
347 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00"),
348 => ("00", "01", "00", "11", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
349 => ("00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00"),
350 => ("00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00"),
351 => ("00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01"),
352 => ("00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01"),
353 => ("00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
354 => ("01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01"),
355 => ("00", "11", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01"),
356 => ("00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01"),
357 => ("00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "01"),
358 => ("01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00"),
359 => ("01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "00"),
360 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
361 => ("00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00"),
362 => ("01", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01"),
363 => ("01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11"),
364 => ("00", "11", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
365 => ("00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "11"),
366 => ("00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "11"),
367 => ("01", "11", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00"),
368 => ("00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
369 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00"),
370 => ("00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01"),
371 => ("01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11"),
372 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "11", "00", "00", "01", "01"),
373 => ("01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01"),
374 => ("00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01"),
375 => ("01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
376 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01"),
377 => ("00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01"),
378 => ("01", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00"),
379 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01"),
380 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "11"),
381 => ("00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00"),
382 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00"),
383 => ("00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00"),
384 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01"),
385 => ("00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01"),
386 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01"),
387 => ("01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
388 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "11", "00", "01", "00"),
389 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01"),
390 => ("00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "11"),
391 => ("01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00"),
392 => ("00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00"),
393 => ("00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "11"),
394 => ("01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01"),
395 => ("01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"),
396 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "01"),
397 => ("01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00"),
398 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00"),
399 => ("00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
400 => ("00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01"),
401 => ("01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11"),
402 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00"),
403 => ("00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00"),
404 => ("00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00"),
405 => ("01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01"),
406 => ("00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11"),
407 => ("01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00"),
408 => ("00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01"),
409 => ("00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "11", "00", "00", "00"),
410 => ("01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00"),
411 => ("01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
412 => ("01", "00", "00", "01", "00", "01", "11", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00"),
413 => ("00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01"),
414 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
415 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01"),
416 => ("00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
417 => ("01", "01", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
418 => ("00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00"),
419 => ("00", "00", "00", "01", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
420 => ("00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
421 => ("01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
422 => ("01", "00", "11", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
423 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01"),
424 => ("00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00"),
425 => ("00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00"),
426 => ("01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01"),
427 => ("01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00"),
428 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "11", "00"),
429 => ("01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
430 => ("00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
431 => ("00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11"),
432 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "11", "01", "01", "01"),
433 => ("00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01"),
434 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
435 => ("00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "11", "00"),
436 => ("00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01"),
437 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00"),
438 => ("01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
439 => ("00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01"),
440 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01"),
441 => ("01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
442 => ("00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00"),
443 => ("00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01"),
444 => ("01", "01", "11", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
445 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11"),
446 => ("00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
447 => ("01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01"),
448 => ("00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00"),
449 => ("00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00"),
450 => ("01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
451 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
452 => ("00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
453 => ("00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01"),
454 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00"),
455 => ("01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00"),
456 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "01"),
457 => ("00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00"),
458 => ("00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "01"),
459 => ("00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
460 => ("01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01"),
461 => ("00", "00", "00", "00", "11", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00"),
462 => ("00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01"),
463 => ("00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01"),
464 => ("00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01"),
465 => ("01", "01", "00", "11", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00"),
466 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11"),
467 => ("00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01"),
468 => ("01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01"),
469 => ("00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
470 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01"),
471 => ("00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
472 => ("01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01"),
473 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
474 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01"),
475 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00"),
476 => ("00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
477 => ("00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00"),
478 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01"),
479 => ("01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01"),
480 => ("01", "11", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01"),
481 => ("01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "11", "00", "01", "01", "01", "01", "00"),
482 => ("01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01"),
483 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "11"),
484 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11"),
485 => ("01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01"),
486 => ("01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
487 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00"),
488 => ("01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11"),
489 => ("01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00"),
490 => ("01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01"),
491 => ("01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00"),
492 => ("00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01"),
493 => ("00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00"),
494 => ("01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
495 => ("01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00"),
496 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01"),
497 => ("00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00"),
498 => ("01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01"),
499 => ("00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "01")),
(
0 => ("01", "01", "11", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
1 => ("01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00"),
2 => ("00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "11", "01", "11", "01", "00", "01", "01", "00", "01"),
3 => ("00", "01", "01", "00", "11", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01"),
4 => ("01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "00"),
5 => ("01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "11", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
6 => ("01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01"),
7 => ("01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
8 => ("00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00"),
9 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00"),
10 => ("00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01"),
11 => ("00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00"),
12 => ("00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
13 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "11", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
14 => ("01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "11", "00", "01", "00", "01", "00"),
15 => ("00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01"),
16 => ("01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01"),
17 => ("01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11"),
18 => ("00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "11", "01", "00", "01", "01", "01"),
19 => ("00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
20 => ("00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01"),
21 => ("01", "01", "00", "11", "01", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
22 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01"),
23 => ("01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01"),
24 => ("00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "11", "00", "00"),
25 => ("00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "11", "11", "01", "01", "00", "00", "01"),
26 => ("00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01"),
27 => ("00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "11", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
28 => ("01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
29 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "11", "00", "01", "00", "01", "11", "01"),
30 => ("00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00"),
31 => ("01", "01", "11", "01", "00", "00", "01", "01", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
32 => ("01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
33 => ("00", "11", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00"),
34 => ("01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01"),
35 => ("01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01"),
36 => ("00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00"),
37 => ("01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01"),
38 => ("00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "11", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01"),
39 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "01", "00", "11", "01"),
40 => ("00", "11", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00"),
41 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "00", "01", "01", "00"),
42 => ("01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01"),
43 => ("00", "01", "11", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
44 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "11", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
45 => ("00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "11", "00", "00"),
46 => ("00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01"),
47 => ("01", "00", "11", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
48 => ("00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01"),
49 => ("01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
50 => ("00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "01"),
51 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "01", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01"),
52 => ("01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01"),
53 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11"),
54 => ("01", "01", "01", "11", "01", "00", "11", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
55 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00"),
56 => ("00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "00"),
57 => ("00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01"),
58 => ("00", "00", "01", "00", "00", "11", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
59 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "11", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00"),
60 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01"),
61 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01", "11", "00"),
62 => ("00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11"),
63 => ("01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01"),
64 => ("01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01"),
65 => ("00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "11", "00", "11"),
66 => ("00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00"),
67 => ("00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "11", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01"),
68 => ("00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00"),
69 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "11", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00"),
70 => ("01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11"),
71 => ("00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00"),
72 => ("01", "01", "01", "11", "11", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00"),
73 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00"),
74 => ("00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00"),
75 => ("01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "01"),
76 => ("01", "00", "01", "11", "00", "11", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
77 => ("00", "11", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01"),
78 => ("00", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01"),
79 => ("01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00"),
80 => ("00", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01"),
81 => ("01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00"),
82 => ("00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11"),
83 => ("01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01"),
84 => ("01", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
85 => ("01", "01", "01", "11", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "00"),
86 => ("00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11"),
87 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00"),
88 => ("01", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01"),
89 => ("01", "00", "01", "00", "01", "11", "00", "11", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
90 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11"),
91 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11"),
92 => ("00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00"),
93 => ("01", "00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01"),
94 => ("01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00"),
95 => ("01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01"),
96 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "11", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01"),
97 => ("01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01"),
98 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "11", "01", "01", "01", "01"),
99 => ("00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "11"),
100 => ("01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
101 => ("01", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01"),
102 => ("00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "00", "00", "01"),
103 => ("00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
104 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00"),
105 => ("01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01"),
106 => ("00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00"),
107 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "11", "11", "01", "00", "00", "00", "01"),
108 => ("01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "11", "01", "00"),
109 => ("00", "00", "00", "00", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00"),
110 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "01", "11", "00", "00", "01"),
111 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01"),
112 => ("00", "01", "11", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11"),
113 => ("01", "01", "01", "01", "01", "01", "01", "11", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01"),
114 => ("01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11"),
115 => ("00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "11", "01"),
116 => ("01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "00", "11"),
117 => ("01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "11", "11", "01", "00", "01", "01", "00", "00", "01", "00"),
118 => ("00", "00", "00", "00", "01", "11", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "01"),
119 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "11", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00"),
120 => ("00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01"),
121 => ("00", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01"),
122 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "11", "01", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
123 => ("01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "11", "00", "00", "01", "00", "00", "00", "01"),
124 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "11", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00"),
125 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "11", "01", "00", "11", "01", "00", "00", "01", "01"),
126 => ("00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
127 => ("00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01"),
128 => ("00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00"),
129 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "11", "01", "11", "01"),
130 => ("00", "00", "00", "00", "11", "11", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
131 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00"),
132 => ("01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00"),
133 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
134 => ("01", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
135 => ("01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
136 => ("00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00"),
137 => ("00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00"),
138 => ("01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "11", "00"),
139 => ("00", "11", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01"),
140 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "11", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00"),
141 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
142 => ("01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01"),
143 => ("00", "01", "11", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
144 => ("01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01"),
145 => ("00", "00", "00", "01", "00", "01", "11", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00"),
146 => ("00", "00", "00", "11", "01", "00", "01", "00", "11", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
147 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "11", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00"),
148 => ("01", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00"),
149 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "11", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01"),
150 => ("01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
151 => ("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "00"),
152 => ("01", "01", "00", "01", "11", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00"),
153 => ("01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00"),
154 => ("00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00"),
155 => ("01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01"),
156 => ("00", "01", "00", "00", "11", "01", "01", "00", "00", "11", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00"),
157 => ("00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01"),
158 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "11", "01", "11", "01", "01", "00", "00", "01", "00"),
159 => ("00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01"),
160 => ("01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "11", "00"),
161 => ("00", "11", "01", "00", "01", "00", "11", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01"),
162 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "00", "11", "11", "01", "01", "00", "01"),
163 => ("01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00"),
164 => ("00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01"),
165 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "00", "01"),
166 => ("01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00"),
167 => ("01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01"),
168 => ("01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
169 => ("00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "00"),
170 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00", "11", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
171 => ("01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "00", "11"),
172 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "01", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
173 => ("00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "00", "11", "01", "01", "00", "11", "01", "00", "01", "01", "01"),
174 => ("00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
175 => ("01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "11", "00", "00", "00", "00"),
176 => ("01", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
177 => ("01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01"),
178 => ("00", "01", "00", "00", "01", "00", "00", "00", "11", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
179 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11"),
180 => ("01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01"),
181 => ("00", "11", "11", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00"),
182 => ("00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01"),
183 => ("00", "00", "01", "00", "01", "00", "11", "00", "11", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
184 => ("01", "01", "01", "00", "01", "01", "11", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
185 => ("00", "00", "11", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00"),
186 => ("01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11"),
187 => ("01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00"),
188 => ("00", "00", "00", "01", "01", "01", "00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00"),
189 => ("00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00"),
190 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "11", "11", "01"),
191 => ("01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00"),
192 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "01", "11", "00"),
193 => ("01", "01", "11", "00", "00", "11", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00"),
194 => ("00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00"),
195 => ("01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00"),
196 => ("00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
197 => ("00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01"),
198 => ("00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "11", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
199 => ("01", "01", "00", "11", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01"),
200 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "11", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11"),
201 => ("01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01"),
202 => ("00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "01"),
203 => ("01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
204 => ("01", "00", "01", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00"),
205 => ("01", "01", "00", "00", "00", "11", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00"),
206 => ("01", "00", "01", "11", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01"),
207 => ("00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "11", "11"),
208 => ("00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00"),
209 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
210 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "00", "11", "00", "11", "01", "00", "01", "00", "00"),
211 => ("00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "11", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01"),
212 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "11", "11", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00"),
213 => ("00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00"),
214 => ("01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "01", "01", "01", "00", "00", "00"),
215 => ("01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
216 => ("01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "01", "11", "01", "00", "01", "00", "00", "01"),
217 => ("00", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
218 => ("00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
219 => ("01", "11", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01"),
220 => ("01", "00", "01", "01", "11", "00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00"),
221 => ("01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11"),
222 => ("00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01"),
223 => ("01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01"),
224 => ("00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00"),
225 => ("00", "00", "00", "11", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00"),
226 => ("01", "01", "01", "01", "00", "01", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01"),
227 => ("01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01"),
228 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01"),
229 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00"),
230 => ("00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01"),
231 => ("00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00"),
232 => ("01", "00", "00", "01", "11", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01"),
233 => ("01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
234 => ("01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "11", "00", "00"),
235 => ("00", "01", "00", "11", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01"),
236 => ("00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01"),
237 => ("00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "11"),
238 => ("01", "00", "00", "00", "00", "01", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00"),
239 => ("01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "00", "11", "00", "00"),
240 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "00"),
241 => ("01", "00", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01"),
242 => ("01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01"),
243 => ("01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01"),
244 => ("00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00", "01", "00", "00", "00", "11"),
245 => ("00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "11", "00", "00", "00"),
246 => ("00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00"),
247 => ("01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "11"),
248 => ("00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00"),
249 => ("00", "00", "11", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
250 => ("00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01"),
251 => ("00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00"),
252 => ("01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "11"),
253 => ("01", "00", "01", "00", "00", "11", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00"),
254 => ("01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00"),
255 => ("00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00"),
256 => ("01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01"),
257 => ("00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "11", "00", "00", "00"),
258 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "11", "00", "01", "00", "01", "00"),
259 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01"),
260 => ("00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "11", "11", "01", "01", "00", "00", "01", "01", "00", "00"),
261 => ("01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "00", "01", "00", "00"),
262 => ("00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "11"),
263 => ("00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
264 => ("00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "11", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
265 => ("00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01"),
266 => ("00", "00", "00", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01"),
267 => ("01", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00"),
268 => ("01", "01", "01", "00", "11", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00"),
269 => ("01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "11", "01", "01"),
270 => ("01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "11", "01", "01", "01", "00", "00", "01"),
271 => ("01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "11"),
272 => ("00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00"),
273 => ("01", "00", "00", "00", "00", "11", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01"),
274 => ("00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
275 => ("00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "11", "01", "00", "00", "01"),
276 => ("01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
277 => ("00", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "11"),
278 => ("00", "01", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01"),
279 => ("00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01"),
280 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00"),
281 => ("00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01"),
282 => ("00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00"),
283 => ("01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "01", "00", "00", "00", "00", "00", "00", "01"),
284 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01"),
285 => ("01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
286 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00"),
287 => ("00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "11"),
288 => ("00", "00", "11", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01"),
289 => ("00", "01", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
290 => ("01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00"),
291 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
292 => ("00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01"),
293 => ("01", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01"),
294 => ("00", "01", "01", "11", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01"),
295 => ("00", "00", "01", "00", "01", "00", "11", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00"),
296 => ("01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "11", "01"),
297 => ("00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01"),
298 => ("00", "00", "11", "00", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
299 => ("00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01"),
300 => ("00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11"),
301 => ("01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00"),
302 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "11", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01"),
303 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01"),
304 => ("01", "01", "01", "01", "01", "01", "01", "11", "11", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
305 => ("00", "11", "01", "00", "00", "00", "11", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01"),
306 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "11", "00", "00", "01", "11", "01", "01", "00", "00", "01"),
307 => ("00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "11", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01"),
308 => ("01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "11", "00", "01", "11", "00", "00"),
309 => ("00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "11", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01"),
310 => ("00", "00", "00", "11", "01", "11", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01"),
311 => ("01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00"),
312 => ("01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "11", "01"),
313 => ("00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00"),
314 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00"),
315 => ("01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00"),
316 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "11", "00", "01", "11", "00", "01", "01", "00", "00"),
317 => ("01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01"),
318 => ("01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "00", "01"),
319 => ("00", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00"),
320 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "11", "01", "01", "11", "01", "01", "00", "00"),
321 => ("00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11"),
322 => ("01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11"),
323 => ("01", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "01"),
324 => ("00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01"),
325 => ("01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "11", "00"),
326 => ("01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01"),
327 => ("01", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00"),
328 => ("01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00"),
329 => ("00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "00"),
330 => ("00", "01", "11", "11", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00"),
331 => ("01", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01"),
332 => ("01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "11", "00", "00", "01"),
333 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "11", "01", "11", "00", "00", "00"),
334 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "11"),
335 => ("01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00"),
336 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00"),
337 => ("00", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00"),
338 => ("01", "11", "00", "01", "11", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
339 => ("00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "00"),
340 => ("00", "00", "11", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00"),
341 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
342 => ("00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00"),
343 => ("00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "00", "00", "00"),
344 => ("01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01"),
345 => ("00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01"),
346 => ("00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01"),
347 => ("01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "01", "01", "01", "01", "00", "00", "01"),
348 => ("01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01"),
349 => ("00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00"),
350 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "11", "00"),
351 => ("00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01"),
352 => ("01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01"),
353 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "00", "11", "00", "00", "00"),
354 => ("00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "01"),
355 => ("01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01"),
356 => ("01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "00", "00", "01", "00", "00", "01", "11", "00"),
357 => ("00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "00", "11", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00"),
358 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01"),
359 => ("01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00"),
360 => ("01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11"),
361 => ("01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "11", "00", "00", "00"),
362 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00"),
363 => ("00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "00"),
364 => ("00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01"),
365 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "11"),
366 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "11"),
367 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "11", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
368 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "11", "01", "01", "01", "00", "00"),
369 => ("01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00"),
370 => ("00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01"),
371 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01"),
372 => ("00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "11", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00"),
373 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00"),
374 => ("01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01"),
375 => ("01", "00", "11", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00"),
376 => ("01", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00"),
377 => ("01", "01", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00"),
378 => ("01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00"),
379 => ("00", "00", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01"),
380 => ("01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
381 => ("01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00"),
382 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "11", "01", "00", "11"),
383 => ("00", "00", "11", "00", "01", "01", "11", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00"),
384 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "11"),
385 => ("01", "00", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01"),
386 => ("00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01"),
387 => ("00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00"),
388 => ("00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01"),
389 => ("00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
390 => ("01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00"),
391 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "11", "11", "01", "11", "00", "00", "00", "00", "00"),
392 => ("00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01"),
393 => ("00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "11"),
394 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "11", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00"),
395 => ("01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01"),
396 => ("00", "01", "01", "01", "11", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01"),
397 => ("00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "11", "01", "11", "00", "00", "00"),
398 => ("00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00"),
399 => ("00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "11", "01", "00", "01"),
400 => ("01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "11", "00"),
401 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "11", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01"),
402 => ("01", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "11", "01", "01"),
403 => ("01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01"),
404 => ("01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00"),
405 => ("00", "11", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
406 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "11", "00", "00", "01", "00"),
407 => ("00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01"),
408 => ("00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00"),
409 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01"),
410 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00"),
411 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "11"),
412 => ("00", "11", "01", "11", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00"),
413 => ("00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "11", "01", "01"),
414 => ("00", "01", "11", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00"),
415 => ("01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01"),
416 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "11", "01", "11"),
417 => ("01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11"),
418 => ("00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01"),
419 => ("00", "00", "11", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01"),
420 => ("01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11"),
421 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "11"),
422 => ("00", "01", "01", "01", "01", "11", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00"),
423 => ("00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "11"),
424 => ("01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01"),
425 => ("01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00"),
426 => ("01", "01", "00", "01", "01", "01", "11", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00"),
427 => ("00", "11", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01"),
428 => ("01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "11", "00"),
429 => ("00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01"),
430 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
431 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00"),
432 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "11", "00", "01"),
433 => ("00", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00"),
434 => ("00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00"),
435 => ("01", "01", "11", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11"),
436 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "00", "11", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
437 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "11", "01"),
438 => ("00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01"),
439 => ("00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01"),
440 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11"),
441 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "11", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
442 => ("00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "11", "00"),
443 => ("00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11"),
444 => ("01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01"),
445 => ("00", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
446 => ("00", "00", "00", "00", "01", "00", "11", "00", "11", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00"),
447 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00"),
448 => ("00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00"),
449 => ("01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00"),
450 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "11", "01", "00", "01"),
451 => ("00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "11"),
452 => ("01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "11", "00", "00", "01"),
453 => ("00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "11", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00"),
454 => ("00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "11", "01", "00", "00"),
455 => ("01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01"),
456 => ("00", "01", "00", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
457 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01"),
458 => ("01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "11", "00"),
459 => ("01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "11", "00"),
460 => ("01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00"),
461 => ("01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "11", "01", "01"),
462 => ("00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "11", "11", "01", "00", "01", "00", "00", "00", "01", "00"),
463 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11"),
464 => ("01", "11", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01"),
465 => ("00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "11", "00", "00", "00"),
466 => ("00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01"),
467 => ("01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "11", "11", "01", "00"),
468 => ("01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00"),
469 => ("01", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
470 => ("01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11"),
471 => ("00", "00", "01", "01", "11", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
472 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01"),
473 => ("00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "11"),
474 => ("00", "00", "11", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01"),
475 => ("00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01"),
476 => ("01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00", "11", "01"),
477 => ("01", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
478 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "11", "01"),
479 => ("00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01"),
480 => ("01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01"),
481 => ("01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01"),
482 => ("00", "11", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00"),
483 => ("00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "01", "11", "01", "00", "00", "00"),
484 => ("01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "00", "01", "00", "01", "01"),
485 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01"),
486 => ("01", "01", "00", "11", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00"),
487 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11"),
488 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
489 => ("00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00"),
490 => ("00", "11", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
491 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
492 => ("00", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01"),
493 => ("01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00"),
494 => ("01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "00", "11", "00", "11", "00"),
495 => ("00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00"),
496 => ("01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "11", "11", "00", "01", "00", "11", "00", "00", "00", "00", "00"),
497 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11"),
498 => ("00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01"),
499 => ("01", "01", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11")),
(
0 => ("00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11"),
1 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "11", "01", "00", "01", "00", "00", "11", "01", "01", "00", "11", "00", "01"),
2 => ("00", "00", "11", "00", "01", "00", "00", "11", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01"),
3 => ("00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "01"),
4 => ("01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "11", "00", "11", "01"),
5 => ("00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "11", "11", "01", "01"),
6 => ("00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "11", "00", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01", "11", "00"),
7 => ("00", "11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"),
8 => ("00", "01", "01", "01", "11", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
9 => ("00", "01", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01"),
10 => ("01", "01", "11", "00", "01", "11", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01"),
11 => ("01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
12 => ("00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "11", "11", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00"),
13 => ("00", "11", "01", "11", "00", "11", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00"),
14 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "01"),
15 => ("01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00"),
16 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "01", "01"),
17 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "11", "11", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00"),
18 => ("00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "11", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00"),
19 => ("00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "01", "00", "11", "00", "00", "11", "01", "00"),
20 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "11", "00", "00", "01", "01", "11", "00", "01", "00", "00", "11"),
21 => ("00", "01", "00", "00", "01", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "11", "11"),
22 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "11", "11", "00", "01", "00", "00", "01", "00", "00"),
23 => ("01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "11", "11", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00"),
24 => ("01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "11", "01", "00"),
25 => ("01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01"),
26 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
27 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00"),
28 => ("00", "01", "00", "01", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "11"),
29 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "11", "01", "11", "01"),
30 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "00", "11"),
31 => ("00", "00", "11", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01"),
32 => ("01", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00"),
33 => ("00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01"),
34 => ("01", "11", "00", "01", "01", "11", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01"),
35 => ("00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00"),
36 => ("00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11"),
37 => ("00", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "11", "11", "00", "01", "00", "00", "00"),
38 => ("01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
39 => ("01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "11", "01", "11", "01", "01", "00", "00", "01"),
40 => ("01", "01", "00", "00", "00", "11", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01"),
41 => ("00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00"),
42 => ("01", "11", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "11", "00"),
43 => ("00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00"),
44 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "11", "00", "11", "11", "01", "00", "00", "01", "00", "00"),
45 => ("01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "11", "00", "00", "00", "00", "00", "01", "01", "11", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
46 => ("01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "11"),
47 => ("01", "11", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01"),
48 => ("01", "11", "00", "00", "00", "11", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01"),
49 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01"),
50 => ("00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01"),
51 => ("00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "11", "11"),
52 => ("00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00"),
53 => ("00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "00", "00", "01"),
54 => ("01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00"),
55 => ("01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11"),
56 => ("01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
57 => ("00", "11", "01", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
58 => ("01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "11", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01"),
59 => ("01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "00", "00"),
60 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "11"),
61 => ("00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01"),
62 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00"),
63 => ("01", "00", "00", "01", "01", "11", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "11", "00", "00"),
64 => ("01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "11", "11", "01", "00", "01", "00", "00", "00", "00", "01"),
65 => ("00", "00", "11", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01"),
66 => ("00", "00", "00", "00", "00", "01", "01", "00", "11", "11", "01", "01", "00", "01", "01", "11", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00"),
67 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "11", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00"),
68 => ("00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "11", "00", "11", "01", "01", "00", "00", "00", "01", "00"),
69 => ("00", "01", "11", "00", "00", "00", "11", "00", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00"),
70 => ("01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "11", "00"),
71 => ("01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01"),
72 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "11", "11", "00"),
73 => ("00", "00", "00", "00", "11", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01"),
74 => ("00", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00"),
75 => ("00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01"),
76 => ("01", "00", "01", "01", "01", "01", "11", "01", "11", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00"),
77 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "11", "00", "00", "00", "01"),
78 => ("00", "11", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01"),
79 => ("00", "00", "00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00"),
80 => ("01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "11", "01", "01", "00", "00", "11", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01"),
81 => ("00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00"),
82 => ("00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01"),
83 => ("01", "00", "01", "01", "01", "00", "01", "11", "01", "11", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01"),
84 => ("01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "11"),
85 => ("00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "11"),
86 => ("00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "11", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00"),
87 => ("00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "11", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
88 => ("01", "01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01"),
89 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "11", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01"),
90 => ("01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00"),
91 => ("01", "11", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01"),
92 => ("01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "11"),
93 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "11", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01"),
94 => ("00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "11", "00"),
95 => ("01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "11", "00"),
96 => ("01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "11", "00", "00", "00", "00"),
97 => ("01", "01", "01", "11", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01"),
98 => ("01", "01", "00", "11", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11"),
99 => ("01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11"),
100 => ("00", "01", "01", "01", "01", "11", "00", "11", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01"),
101 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "11", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00"),
102 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "01", "11", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00"),
103 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "11", "01"),
104 => ("00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00"),
105 => ("01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "11", "01", "00", "00", "01", "01", "11", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
106 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "11", "00", "00", "11", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01"),
107 => ("01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11", "01", "01", "01", "01", "01", "00", "11", "11", "00", "00", "00"),
108 => ("00", "11", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "11"),
109 => ("00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "11", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00"),
110 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00", "00"),
111 => ("00", "11", "11", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01"),
112 => ("00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01"),
113 => ("01", "11", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01"),
114 => ("01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01"),
115 => ("01", "11", "00", "00", "00", "01", "11", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01"),
116 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "11", "01", "00", "01", "01", "01", "11", "01", "01", "01", "11", "00", "00"),
117 => ("01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "11", "11", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01"),
118 => ("01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01"),
119 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00"),
120 => ("01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01"),
121 => ("00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
122 => ("01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11"),
123 => ("00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01"),
124 => ("00", "00", "11", "01", "01", "01", "00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00"),
125 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "11", "01", "01", "01", "11", "01"),
126 => ("00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "01", "01", "01", "11", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
127 => ("01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00"),
128 => ("00", "11", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "11", "00", "01"),
129 => ("00", "11", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01"),
130 => ("00", "01", "11", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11"),
131 => ("00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "11", "01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01"),
132 => ("01", "00", "01", "00", "01", "11", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00"),
133 => ("01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "11", "11", "00", "01"),
134 => ("00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01"),
135 => ("01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00"),
136 => ("01", "00", "00", "01", "01", "11", "11", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00"),
137 => ("00", "00", "00", "11", "01", "00", "00", "00", "11", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01"),
138 => ("01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "01"),
139 => ("00", "11", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00"),
140 => ("00", "00", "01", "01", "11", "01", "00", "11", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01"),
141 => ("00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "11", "01", "00", "01"),
142 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "01"),
143 => ("01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "11", "00", "00", "01", "01"),
144 => ("01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
145 => ("00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "00", "11", "00", "01", "01", "11", "01", "01", "01", "01", "11", "01"),
146 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "01"),
147 => ("00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "11", "01", "11", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01"),
148 => ("01", "01", "11", "01", "01", "01", "11", "00", "11", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
149 => ("00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00"),
150 => ("01", "00", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11"),
151 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "00", "11", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11"),
152 => ("01", "11", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00"),
153 => ("00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "11", "00", "11"),
154 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "11", "00"),
155 => ("01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "00", "00", "01", "11", "00", "11", "00", "00", "01", "00"),
156 => ("00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
157 => ("00", "11", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "00", "11", "01", "00", "01"),
158 => ("00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "00", "11", "11", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01"),
159 => ("00", "01", "11", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01"),
160 => ("00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00"),
161 => ("01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01"),
162 => ("01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "11", "01"),
163 => ("01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "11", "01", "00", "11", "00", "00"),
164 => ("01", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "11", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00"),
165 => ("01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "11", "11", "01", "01", "01", "00", "01", "01", "11", "00"),
166 => ("00", "00", "01", "11", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "00"),
167 => ("01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "11", "11", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01"),
168 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "11", "00", "11", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
169 => ("01", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "11", "00", "11", "00", "00", "01"),
170 => ("00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "11", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11"),
171 => ("00", "01", "01", "11", "11", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00"),
172 => ("01", "00", "00", "00", "00", "11", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00"),
173 => ("01", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "11", "00", "11", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
174 => ("00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "11", "11", "00", "11"),
175 => ("00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00"),
176 => ("01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "11", "01", "00", "01", "00", "00", "00"),
177 => ("00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "11", "00"),
178 => ("01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "11", "01", "01", "00"),
179 => ("01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01"),
180 => ("01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "00", "01", "00", "11", "11", "01", "00", "00", "01"),
181 => ("01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00"),
182 => ("01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "11", "01", "11", "00", "00", "00", "01", "00", "01", "00", "11", "00"),
183 => ("00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00"),
184 => ("00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00"),
185 => ("00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "00"),
186 => ("01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "11", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "00"),
187 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "11", "01", "01", "11", "00", "01"),
188 => ("00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "11", "11", "00", "00", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
189 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "01", "11", "01", "01"),
190 => ("00", "11", "00", "00", "01", "11", "11", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
191 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "11", "01", "00", "00", "00"),
192 => ("01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
193 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "11", "11", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
194 => ("00", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "01", "00"),
195 => ("00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "00", "01", "01", "01", "01"),
196 => ("01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00"),
197 => ("01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01"),
198 => ("01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "11", "01", "11", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00"),
199 => ("00", "01", "01", "01", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00"),
200 => ("00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "11", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00"),
201 => ("01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11"),
202 => ("01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "11", "11", "00", "00"),
203 => ("00", "00", "11", "11", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00"),
204 => ("00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "11", "01"),
205 => ("01", "11", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00"),
206 => ("01", "11", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11"),
207 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "11", "00", "00"),
208 => ("00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
209 => ("00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01"),
210 => ("01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00"),
211 => ("01", "00", "01", "01", "00", "11", "11", "00", "01", "01", "01", "11", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
212 => ("01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "11", "01", "11", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01"),
213 => ("00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01"),
214 => ("00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
215 => ("00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00"),
216 => ("00", "01", "00", "11", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "11", "01", "00"),
217 => ("00", "01", "01", "01", "01", "01", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01"),
218 => ("01", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "11", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00"),
219 => ("01", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01"),
220 => ("01", "00", "11", "01", "01", "11", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00"),
221 => ("01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01"),
222 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "11", "01", "01"),
223 => ("01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01"),
224 => ("00", "00", "01", "01", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01"),
225 => ("01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00"),
226 => ("00", "11", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "11", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
227 => ("01", "00", "00", "11", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00"),
228 => ("00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01"),
229 => ("00", "11", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "11", "01"),
230 => ("00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01"),
231 => ("01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "00", "11", "11", "11", "01", "00", "00", "00", "01", "01", "01", "00"),
232 => ("00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "00", "01", "00"),
233 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00"),
234 => ("00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "11", "11", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00"),
235 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "11"),
236 => ("01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "11", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01"),
237 => ("00", "11", "01", "00", "00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01"),
238 => ("01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "11", "01"),
239 => ("00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00"),
240 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "11", "00", "00", "01", "11", "01", "01", "00", "01", "11", "01", "00", "01", "01"),
241 => ("00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "11", "11", "00", "11", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00"),
242 => ("00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "11", "00", "00", "00"),
243 => ("00", "11", "00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01"),
244 => ("01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "11", "01", "01"),
245 => ("00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "11", "00"),
246 => ("00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00"),
247 => ("00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
248 => ("01", "00", "01", "11", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01"),
249 => ("01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "01", "11", "00"),
250 => ("01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "11", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
251 => ("00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "11", "00", "01", "01", "11", "01", "00", "00", "00", "01"),
252 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "11", "01"),
253 => ("00", "00", "01", "11", "11", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01"),
254 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "11", "01", "11", "01", "01"),
255 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "11", "01", "01", "00", "00"),
256 => ("01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
257 => ("00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11"),
258 => ("01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "11"),
259 => ("00", "00", "01", "11", "00", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01"),
260 => ("00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "11", "00", "11", "00"),
261 => ("01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "01", "01", "11"),
262 => ("00", "00", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00"),
263 => ("00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "11", "01"),
264 => ("01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00"),
265 => ("00", "11", "00", "11", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00"),
266 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "11", "00", "00", "00", "11", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01"),
267 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "11", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00"),
268 => ("01", "01", "00", "00", "11", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "11"),
269 => ("00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "11", "00", "01", "11", "00", "01", "01", "00", "00", "00", "11"),
270 => ("01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00"),
271 => ("01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "11", "01", "01", "01"),
272 => ("01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01"),
273 => ("01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00"),
274 => ("01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01"),
275 => ("00", "01", "01", "01", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01"),
276 => ("00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "11", "00", "11", "00", "01"),
277 => ("01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "00"),
278 => ("00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "11", "00", "00", "11", "01", "00", "01", "00", "00", "01"),
279 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "11"),
280 => ("01", "11", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00"),
281 => ("00", "01", "01", "01", "11", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01"),
282 => ("00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "11", "00", "01", "00"),
283 => ("00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01"),
284 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "11", "11", "01", "00", "00"),
285 => ("00", "00", "11", "01", "00", "01", "11", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01"),
286 => ("00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "11", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01"),
287 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "11", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00"),
288 => ("01", "11", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00"),
289 => ("00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "11", "00", "00"),
290 => ("00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01"),
291 => ("00", "01", "01", "01", "01", "01", "00", "11", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "00"),
292 => ("00", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01"),
293 => ("00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "11", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00"),
294 => ("01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "11", "01", "00"),
295 => ("00", "01", "01", "11", "01", "00", "00", "01", "00", "11", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00"),
296 => ("00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00", "01", "11", "00", "11", "01", "00", "01", "01", "00"),
297 => ("01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "11", "11", "01", "01", "01"),
298 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "11", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "11", "00"),
299 => ("00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "01"),
300 => ("01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00"),
301 => ("00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00"),
302 => ("01", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11"),
303 => ("01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01"),
304 => ("01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "11", "01", "11", "01", "00", "01"),
305 => ("01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "11", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01"),
306 => ("00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01"),
307 => ("00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11"),
308 => ("00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00"),
309 => ("00", "00", "01", "01", "11", "00", "11", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00"),
310 => ("00", "00", "00", "11", "11", "01", "11", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01"),
311 => ("00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "11", "01", "01"),
312 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "11", "01"),
313 => ("01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "11"),
314 => ("01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01"),
315 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "01", "11", "00", "11", "00", "01"),
316 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
317 => ("00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "11", "00", "00", "11", "00", "01", "00"),
318 => ("01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "11", "00", "00", "01", "00", "00", "00"),
319 => ("00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00"),
320 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "11", "11", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00"),
321 => ("01", "01", "01", "00", "01", "11", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00"),
322 => ("01", "00", "11", "00", "11", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00"),
323 => ("01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "11", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00"),
324 => ("01", "01", "00", "11", "00", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
325 => ("01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "11", "01"),
326 => ("01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "00", "00"),
327 => ("00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "11", "00", "00"),
328 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "11"),
329 => ("01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "01", "11", "01", "00", "01", "11", "01"),
330 => ("01", "11", "01", "00", "00", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00"),
331 => ("00", "00", "00", "00", "00", "01", "00", "11", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00"),
332 => ("01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "11", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00"),
333 => ("01", "01", "00", "01", "01", "00", "00", "11", "00", "11", "11", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00"),
334 => ("01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00"),
335 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "11", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00"),
336 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "11", "11", "01", "11", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00"),
337 => ("01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00"),
338 => ("01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01"),
339 => ("01", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "00", "00", "00", "00"),
340 => ("00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "11", "11", "01", "00", "01", "00", "00", "00", "00", "00"),
341 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01"),
342 => ("01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "11", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00"),
343 => ("00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "00", "01", "11", "00", "00", "01", "01"),
344 => ("01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "11", "11", "01", "11", "01"),
345 => ("00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11"),
346 => ("00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11"),
347 => ("00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00"),
348 => ("01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "11"),
349 => ("00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "01"),
350 => ("01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "00", "11", "01", "11", "00"),
351 => ("01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "11", "11", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01"),
352 => ("01", "11", "00", "00", "01", "11", "01", "00", "00", "01", "01", "11", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
353 => ("01", "00", "00", "01", "11", "00", "01", "00", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00"),
354 => ("00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
355 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "11", "11"),
356 => ("00", "00", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "01", "00", "00", "00"),
357 => ("00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "11", "01", "01"),
358 => ("00", "00", "01", "00", "11", "11", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01"),
359 => ("00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01"),
360 => ("00", "11", "00", "00", "00", "11", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01"),
361 => ("00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "11", "01", "01", "01"),
362 => ("01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01"),
363 => ("01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "11", "01", "01", "00", "11", "11", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
364 => ("01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00"),
365 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "01"),
366 => ("01", "00", "11", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "11", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00"),
367 => ("00", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "11", "01", "01", "11", "01", "11"),
368 => ("00", "11", "01", "01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00"),
369 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "00", "01", "01"),
370 => ("00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "11", "01", "01", "01", "01", "11", "01", "11"),
371 => ("00", "00", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11"),
372 => ("00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00"),
373 => ("00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00"),
374 => ("00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "11", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01"),
375 => ("00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "11", "01", "01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00"),
376 => ("00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01"),
377 => ("01", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "00", "01", "00", "01", "11", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00"),
378 => ("01", "01", "00", "00", "01", "01", "11", "11", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01"),
379 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "11", "01", "11", "11", "01", "00", "01", "00", "00", "01", "01"),
380 => ("00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00"),
381 => ("01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "11", "00", "01", "00", "00", "01", "01", "01", "00", "11"),
382 => ("00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00"),
383 => ("01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "11", "01", "00", "01", "00", "01", "11", "01", "00"),
384 => ("00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00"),
385 => ("01", "00", "00", "11", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00"),
386 => ("00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11"),
387 => ("00", "11", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00"),
388 => ("01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "11", "01", "00", "00", "01", "00"),
389 => ("00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "11", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "00", "01"),
390 => ("01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "00"),
391 => ("00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "01", "11", "11"),
392 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "11", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01"),
393 => ("01", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00"),
394 => ("00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01"),
395 => ("01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "00", "01"),
396 => ("01", "00", "11", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01"),
397 => ("00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00"),
398 => ("00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "01", "00", "01", "11", "00"),
399 => ("01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "11", "01", "00", "00", "00", "11", "01"),
400 => ("00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01"),
401 => ("00", "01", "01", "01", "11", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00"),
402 => ("01", "01", "01", "00", "11", "11", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01"),
403 => ("01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "01", "00"),
404 => ("00", "01", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00"),
405 => ("00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01"),
406 => ("00", "11", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "11", "00", "00"),
407 => ("00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00"),
408 => ("01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01"),
409 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "11", "01", "01", "00", "00", "11", "01"),
410 => ("00", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "11", "00", "00", "11", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00"),
411 => ("01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01"),
412 => ("01", "11", "01", "11", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00"),
413 => ("00", "11", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "11", "01", "01", "01"),
414 => ("01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "11", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00"),
415 => ("01", "01", "01", "00", "11", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11"),
416 => ("01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00"),
417 => ("00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "11", "00", "01", "00", "11"),
418 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "11", "00", "00", "00", "01", "01", "01", "11", "11", "00", "01", "01", "00", "00"),
419 => ("00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "01", "00"),
420 => ("00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "11", "01", "00", "01", "01", "11", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00"),
421 => ("01", "01", "01", "11", "00", "00", "01", "11", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01"),
422 => ("00", "00", "11", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "00"),
423 => ("00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01"),
424 => ("00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00"),
425 => ("01", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "11"),
426 => ("01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00"),
427 => ("00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01"),
428 => ("01", "01", "01", "00", "11", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00"),
429 => ("01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "11", "11", "01", "11", "01", "01", "01", "00", "00"),
430 => ("01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "11", "11", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
431 => ("01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "11", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "00", "00"),
432 => ("01", "00", "01", "11", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00"),
433 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
434 => ("00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "11", "01", "11", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01"),
435 => ("00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01"),
436 => ("00", "11", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01"),
437 => ("01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "11", "00", "11", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00"),
438 => ("01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00", "11", "01"),
439 => ("00", "00", "00", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01"),
440 => ("00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01"),
441 => ("01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "01"),
442 => ("01", "00", "00", "00", "01", "01", "11", "00", "00", "11", "01", "00", "01", "11", "00", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01"),
443 => ("01", "00", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00"),
444 => ("01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00"),
445 => ("01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "11", "00", "01", "11", "00", "01", "00", "11", "01"),
446 => ("01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "00", "00"),
447 => ("01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00"),
448 => ("00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "11", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "00"),
449 => ("00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "11", "00", "01", "01", "00", "00", "01"),
450 => ("01", "01", "00", "11", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "11", "01", "00", "00", "01"),
451 => ("01", "00", "00", "00", "11", "11", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00"),
452 => ("00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01"),
453 => ("01", "11", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "01", "11", "00", "00", "11", "01", "01"),
454 => ("00", "01", "01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00"),
455 => ("00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "11", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00"),
456 => ("00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "11", "00", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "00"),
457 => ("00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "11", "01"),
458 => ("01", "11", "01", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00"),
459 => ("01", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "01", "11", "01"),
460 => ("01", "11", "00", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00"),
461 => ("01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11", "01", "01", "00", "11", "00", "01", "01", "11", "00", "01", "01", "00"),
462 => ("00", "01", "01", "01", "01", "01", "01", "01", "11", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "01", "00", "00", "01", "00", "01"),
463 => ("00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "11"),
464 => ("00", "01", "11", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "01", "00", "11", "00", "01"),
465 => ("01", "01", "01", "11", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00"),
466 => ("00", "01", "11", "00", "11", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
467 => ("01", "01", "11", "01", "01", "00", "00", "11", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "01"),
468 => ("00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01"),
469 => ("00", "00", "00", "00", "01", "01", "11", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "11", "00"),
470 => ("01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "11"),
471 => ("01", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00"),
472 => ("00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "11", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00"),
473 => ("00", "01", "01", "11", "00", "01", "01", "01", "01", "11", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01"),
474 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00"),
475 => ("01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01"),
476 => ("00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "11", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01"),
477 => ("00", "01", "00", "00", "01", "00", "11", "11", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01"),
478 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "00", "11", "11"),
479 => ("00", "11", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01"),
480 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "11", "01", "11", "11", "01", "00", "00", "00", "01", "01"),
481 => ("01", "11", "11", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01"),
482 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "11", "00"),
483 => ("00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "11", "00", "00", "11"),
484 => ("01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "11"),
485 => ("01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11"),
486 => ("00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "11", "01", "11", "01", "00", "00"),
487 => ("00", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "11", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00"),
488 => ("01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "11", "01", "11", "01", "01", "01", "01"),
489 => ("01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11"),
490 => ("01", "00", "00", "00", "11", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "11", "01", "01", "00", "01"),
491 => ("00", "11", "01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
492 => ("00", "00", "11", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "11", "01", "01", "01"),
493 => ("00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "11", "01", "01", "01"),
494 => ("01", "01", "01", "00", "11", "01", "11", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00"),
495 => ("01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01"),
496 => ("01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "11", "11", "01", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
497 => ("01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "11", "00", "01", "01", "00", "01", "01", "01"),
498 => ("00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00"),
499 => ("00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00")),
(
0 => ("01", "01", "00", "11", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "11", "01", "11", "01", "00", "00", "00"),
1 => ("00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01"),
2 => ("01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00"),
3 => ("00", "00", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00"),
4 => ("01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "00", "00", "00", "00", "11", "01", "00"),
5 => ("01", "00", "01", "11", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "11", "01", "00", "11"),
6 => ("01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00", "11", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "11"),
7 => ("00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "11", "01"),
8 => ("01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "11", "11", "00", "00", "01", "11", "01", "00", "00"),
9 => ("00", "11", "00", "11", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "11", "01", "00", "00", "00", "00"),
10 => ("01", "11", "00", "01", "11", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00"),
11 => ("00", "01", "11", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01"),
12 => ("00", "01", "01", "01", "11", "00", "00", "00", "11", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "11", "01", "01", "01", "01"),
13 => ("00", "00", "11", "00", "00", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00"),
14 => ("01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
15 => ("00", "00", "11", "00", "00", "01", "00", "11", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01"),
16 => ("00", "00", "00", "11", "00", "00", "11", "00", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "11", "00", "00"),
17 => ("00", "11", "11", "01", "11", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00"),
18 => ("01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "11", "00", "01", "11"),
19 => ("00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "11", "11", "01", "00", "01", "01", "01", "01", "11", "01", "00", "11", "01", "00", "00"),
20 => ("00", "01", "11", "00", "01", "00", "01", "11", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "11"),
21 => ("00", "01", "01", "01", "01", "11", "11", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "11"),
22 => ("00", "01", "00", "11", "00", "00", "00", "11", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01"),
23 => ("00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "11", "11", "01", "00", "00", "01", "01"),
24 => ("00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "01", "11", "11", "11", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01"),
25 => ("01", "11", "00", "00", "11", "11", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
26 => ("00", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "11", "01", "00", "00", "00"),
27 => ("01", "11", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01"),
28 => ("00", "00", "01", "11", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11"),
29 => ("01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "11", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "11"),
30 => ("01", "11", "01", "11", "01", "01", "01", "01", "11", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00"),
31 => ("00", "00", "00", "01", "00", "11", "00", "01", "01", "11", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00"),
32 => ("01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "11", "01", "11", "01", "00"),
33 => ("01", "01", "01", "00", "11", "11", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "00", "00", "01"),
34 => ("00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "11", "01", "00", "11", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00"),
35 => ("01", "01", "01", "11", "01", "00", "00", "11", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "00", "01"),
36 => ("00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "11"),
37 => ("01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "11", "00", "00", "01", "01", "11", "01", "01", "01", "00", "11", "00", "01", "00", "11", "01", "00", "00", "01"),
38 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "11", "00", "00", "11", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "11", "11"),
39 => ("01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "11", "01", "11", "11", "00"),
40 => ("00", "01", "01", "11", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "11", "01", "01", "01", "01", "01"),
41 => ("00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11"),
42 => ("00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "11", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00", "00"),
43 => ("00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "11", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01"),
44 => ("01", "00", "01", "01", "01", "00", "11", "11", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "11", "01"),
45 => ("00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01"),
46 => ("00", "00", "00", "00", "11", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "11", "11", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
47 => ("01", "01", "01", "01", "00", "11", "00", "11", "01", "11", "11", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
48 => ("01", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "11"),
49 => ("00", "01", "01", "00", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00"),
50 => ("00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "11", "00", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01"),
51 => ("00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01"),
52 => ("00", "01", "11", "01", "11", "11", "01", "00", "11", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01"),
53 => ("01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00"),
54 => ("01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "11", "11", "11", "00", "00", "00", "00", "01"),
55 => ("00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "11", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01"),
56 => ("00", "11", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "11", "00", "00", "01"),
57 => ("01", "11", "11", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00"),
58 => ("00", "11", "01", "00", "11", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01"),
59 => ("00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "11", "11", "01", "01", "00", "01", "11", "01", "00", "00"),
60 => ("01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00"),
61 => ("00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "11", "00", "01", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00"),
62 => ("01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "11", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "11"),
63 => ("00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "01", "11", "00", "01", "00", "00", "01", "11", "01"),
64 => ("01", "00", "00", "00", "11", "00", "11", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "11", "00"),
65 => ("01", "11", "00", "01", "00", "11", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01"),
66 => ("01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "11", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
67 => ("00", "00", "01", "01", "11", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "00"),
68 => ("01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "11", "11", "01"),
69 => ("01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "11", "11", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "01", "11"),
70 => ("00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00"),
71 => ("00", "00", "11", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "11", "01"),
72 => ("00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00"),
73 => ("00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "11", "00", "00"),
74 => ("01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "11", "01", "01", "11", "11", "01", "01", "00", "00", "00", "11", "00", "00"),
75 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "11", "00", "11", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00"),
76 => ("00", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "11", "00", "01", "01", "00", "01", "00", "01", "11", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01"),
77 => ("00", "01", "11", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "11", "00", "01", "01", "01", "11", "01"),
78 => ("01", "00", "11", "11", "01", "00", "01", "01", "11", "01", "11", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01"),
79 => ("00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "01", "11", "01", "00", "00", "11", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00"),
80 => ("01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "11", "01", "11", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00"),
81 => ("00", "01", "11", "01", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "11", "11", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01"),
82 => ("00", "01", "01", "01", "11", "00", "11", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "01", "01"),
83 => ("01", "01", "11", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00"),
84 => ("00", "11", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "01", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01"),
85 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "11", "00", "00", "01", "11", "00", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00"),
86 => ("00", "00", "00", "01", "00", "01", "11", "01", "00", "11", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00"),
87 => ("00", "00", "01", "00", "11", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "11", "01", "11", "00", "00", "00", "01", "01", "01", "00"),
88 => ("00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "11", "00", "11", "01"),
89 => ("01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "00", "01", "00"),
90 => ("00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "11", "11", "11", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01"),
91 => ("01", "01", "00", "00", "00", "11", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "11"),
92 => ("00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "00", "01", "01", "11"),
93 => ("00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "11", "01", "00", "01", "00", "01", "00", "01", "11", "11", "01", "00"),
94 => ("01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11"),
95 => ("01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00", "11", "11", "11", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01"),
96 => ("01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "11", "11", "00", "01", "00"),
97 => ("00", "00", "00", "00", "00", "11", "11", "11", "00", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00"),
98 => ("00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00", "11", "00", "00", "00", "00", "01", "11", "00", "01"),
99 => ("00", "00", "00", "01", "01", "01", "11", "11", "01", "01", "01", "00", "00", "01", "00", "11", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
100 => ("00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "00", "11"),
101 => ("00", "00", "00", "01", "11", "11", "01", "01", "00", "01", "01", "11", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "01", "00", "01"),
102 => ("00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00", "00", "00"),
103 => ("01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11", "00", "01", "00", "00"),
104 => ("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "11", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00"),
105 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01", "01", "11", "11", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01"),
106 => ("00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "11", "00", "01", "01", "00", "11"),
107 => ("00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "11", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "11", "00", "00"),
108 => ("01", "11", "11", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00"),
109 => ("00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00"),
110 => ("01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "00", "11", "00", "00"),
111 => ("01", "00", "00", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "11", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
112 => ("00", "11", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "00", "11", "01"),
113 => ("00", "11", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00"),
114 => ("00", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01"),
115 => ("01", "11", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "11", "01", "00", "00", "11", "00", "00", "01"),
116 => ("01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "11", "01", "00", "00", "11", "01", "00", "11", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01"),
117 => ("00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
118 => ("00", "01", "11", "00", "00", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "11", "00"),
119 => ("00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "11"),
120 => ("01", "11", "01", "11", "00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00"),
121 => ("01", "00", "11", "00", "00", "00", "01", "01", "11", "11", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00"),
122 => ("01", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "11", "01", "01", "11", "00"),
123 => ("00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "11", "00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
124 => ("01", "00", "01", "00", "01", "11", "01", "01", "11", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00"),
125 => ("00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "11", "01", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "01"),
126 => ("01", "01", "00", "00", "11", "00", "01", "01", "01", "11", "01", "01", "01", "11", "00", "11", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01"),
127 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "11", "11", "00", "11", "00", "00", "01", "01", "11", "01", "00", "01"),
128 => ("01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00"),
129 => ("00", "00", "00", "00", "11", "01", "00", "01", "11", "01", "11", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00"),
130 => ("00", "01", "00", "00", "11", "00", "01", "00", "00", "11", "01", "01", "11", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01"),
131 => ("01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "11", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "11", "11", "00"),
132 => ("01", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11"),
133 => ("00", "00", "01", "01", "00", "11", "00", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00"),
134 => ("01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "11", "01", "11", "01", "00", "01", "00", "00", "01", "01"),
135 => ("01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "01"),
136 => ("01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "11", "11", "11", "00", "00", "00", "01"),
137 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "11", "00", "01", "11", "01", "11", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01"),
138 => ("01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01"),
139 => ("00", "00", "00", "01", "11", "00", "00", "00", "11", "11", "01", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01"),
140 => ("01", "00", "01", "01", "00", "01", "11", "11", "11", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01"),
141 => ("01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "11", "11", "01", "01", "01", "01", "11", "00"),
142 => ("01", "01", "11", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "11", "00", "11", "00", "00", "01", "01", "01"),
143 => ("01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "11", "01"),
144 => ("01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01"),
145 => ("00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00"),
146 => ("00", "11", "00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00"),
147 => ("00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "00", "11", "11", "00", "01", "00", "01", "11", "00"),
148 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "11", "01", "11", "00", "01", "01"),
149 => ("01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "11", "11", "01", "00", "01", "01", "00", "00", "00", "11"),
150 => ("00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "11", "00", "11", "01", "00", "00", "01", "01", "00", "01", "11"),
151 => ("01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01"),
152 => ("01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "11", "11", "01", "00"),
153 => ("00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "01", "11", "00", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01"),
154 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "11", "11", "00", "00", "11", "00", "00", "00", "00"),
155 => ("01", "00", "11", "00", "00", "00", "11", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01"),
156 => ("01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "11", "01", "01", "11", "00", "01", "01", "11", "00", "11", "00", "01", "01", "01", "00", "01", "00"),
157 => ("01", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00"),
158 => ("01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "11", "00", "01"),
159 => ("01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00"),
160 => ("00", "00", "00", "11", "00", "11", "00", "11", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00"),
161 => ("00", "00", "00", "11", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01"),
162 => ("01", "00", "00", "01", "00", "01", "00", "11", "11", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01"),
163 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "11", "00", "00", "00", "01", "00", "01", "01", "11", "11", "00", "01", "00"),
164 => ("00", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00"),
165 => ("01", "00", "01", "11", "00", "11", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "00", "11", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00"),
166 => ("01", "11", "01", "00", "11", "00", "01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "11", "01"),
167 => ("01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00"),
168 => ("00", "01", "00", "00", "01", "11", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00"),
169 => ("01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "11", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00"),
170 => ("00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "11", "11", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00"),
171 => ("01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "11", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "11", "00"),
172 => ("01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "00", "11", "01"),
173 => ("01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "11", "00", "11", "00"),
174 => ("00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "00"),
175 => ("01", "00", "11", "01", "01", "01", "01", "01", "01", "11", "01", "01", "11", "00", "01", "11", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01"),
176 => ("01", "01", "11", "00", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01"),
177 => ("01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "11", "00", "00", "00", "11", "11", "01", "00", "01", "00", "00"),
178 => ("00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "00", "11", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01"),
179 => ("01", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "01", "00", "01", "11", "11", "01", "01", "00", "01", "01", "00", "01"),
180 => ("01", "01", "01", "11", "00", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "00", "00", "00"),
181 => ("01", "01", "01", "01", "01", "11", "01", "00", "11", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01"),
182 => ("00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "11", "00"),
183 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "11", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "01", "11", "01"),
184 => ("01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "11", "01", "01", "00", "11", "00", "11", "00", "01", "01"),
185 => ("00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "11", "00", "00", "01", "11", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01"),
186 => ("00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "11"),
187 => ("00", "00", "01", "11", "11", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "01"),
188 => ("01", "00", "00", "00", "11", "11", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01"),
189 => ("00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "11", "01", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00"),
190 => ("01", "01", "01", "01", "11", "00", "11", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
191 => ("01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "11", "01", "00", "01", "00", "11", "01", "00", "00", "00"),
192 => ("01", "00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "11", "00", "00"),
193 => ("01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "11", "00", "11", "00"),
194 => ("01", "11", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "11", "01", "11", "01", "00", "00", "00", "00", "00", "00"),
195 => ("00", "11", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00"),
196 => ("01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00"),
197 => ("00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "11", "01", "00"),
198 => ("00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "11", "11", "11", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00"),
199 => ("01", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "01", "01", "11", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "00"),
200 => ("01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "01", "00", "01"),
201 => ("00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "11", "00", "01", "11", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00"),
202 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "11", "01", "11", "00", "01"),
203 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "11", "00", "01", "01", "11", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01"),
204 => ("00", "00", "01", "01", "01", "00", "00", "11", "11", "00", "01", "00", "11", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01"),
205 => ("00", "01", "00", "00", "00", "11", "11", "01", "00", "01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00"),
206 => ("01", "00", "11", "00", "00", "00", "11", "01", "00", "00", "11", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01"),
207 => ("00", "00", "00", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01"),
208 => ("00", "00", "11", "00", "01", "00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00"),
209 => ("01", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "11", "00", "01", "00", "01", "11", "00", "00", "01", "00", "11", "00", "01", "01"),
210 => ("01", "00", "11", "00", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01"),
211 => ("01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "11", "01", "01", "11", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
212 => ("01", "00", "01", "01", "00", "00", "01", "00", "11", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "00", "00"),
213 => ("01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "00", "00", "01", "01", "11", "11", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00"),
214 => ("01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "00", "00", "11", "01", "11", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00"),
215 => ("01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00", "00", "00", "00", "01", "11", "11", "00", "00", "01"),
216 => ("01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01"),
217 => ("01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "11", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "01", "01", "00", "01", "00"),
218 => ("00", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "11", "00", "11", "00", "01", "01", "00", "01", "11", "00", "00", "01"),
219 => ("01", "00", "00", "11", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01"),
220 => ("01", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00"),
221 => ("01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "11", "11", "00", "01", "01"),
222 => ("00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "11", "11", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00"),
223 => ("01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "11", "00", "00", "11", "00", "01", "01", "11", "00", "11", "01", "01", "00"),
224 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "11", "00", "01", "00", "01", "11", "01", "11", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00"),
225 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "01", "11", "01", "00", "11", "01", "00", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "00", "00"),
226 => ("01", "00", "00", "11", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01"),
227 => ("01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "00", "11", "11", "00", "11", "01", "11", "01", "00", "00"),
228 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "11", "00", "11", "01", "01", "01", "00", "01", "11", "11", "01", "00", "00"),
229 => ("01", "01", "11", "01", "00", "11", "01", "01", "00", "00", "11", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01"),
230 => ("00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "01", "11", "00", "01", "01"),
231 => ("01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "11", "00", "11", "00", "01", "11", "01", "00", "01", "00"),
232 => ("01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "11", "01", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00"),
233 => ("00", "00", "01", "00", "00", "00", "11", "01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11"),
234 => ("01", "11", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "11", "11", "01", "00", "00", "00", "01"),
235 => ("00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "11", "11", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01"),
236 => ("01", "00", "01", "00", "11", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00"),
237 => ("01", "01", "11", "01", "00", "00", "11", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "01"),
238 => ("01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "11", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "11", "00"),
239 => ("01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "00", "00"),
240 => ("00", "11", "01", "11", "01", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01"),
241 => ("00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "11", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01"),
242 => ("00", "01", "01", "00", "01", "01", "01", "00", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00"),
243 => ("01", "11", "00", "01", "11", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "01", "11", "01", "01"),
244 => ("00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "11", "11", "01", "00", "01", "01", "00", "00"),
245 => ("01", "00", "00", "01", "01", "00", "00", "11", "00", "11", "01", "11", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00"),
246 => ("00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "11", "00", "11", "01", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01"),
247 => ("01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "00", "01"),
248 => ("00", "01", "00", "11", "01", "11", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "11", "00"),
249 => ("00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "11", "11", "00", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00"),
250 => ("00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "11", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01"),
251 => ("00", "01", "01", "01", "11", "00", "00", "11", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00"),
252 => ("01", "11", "00", "11", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "11", "00", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01"),
253 => ("01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "11", "00", "00"),
254 => ("01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "11", "00", "01", "11", "01", "00", "01"),
255 => ("00", "01", "11", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00"),
256 => ("00", "01", "11", "01", "01", "11", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "11"),
257 => ("00", "00", "11", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "11", "00", "01", "00", "00", "11", "01", "01", "01", "01"),
258 => ("01", "01", "01", "00", "00", "01", "11", "00", "01", "00", "11", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01"),
259 => ("00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "11", "00", "00", "00", "11", "00", "00", "00", "11"),
260 => ("01", "01", "11", "11", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "11", "01", "00", "01", "01", "01", "00", "00", "11", "01"),
261 => ("00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "11", "11", "01", "01", "01", "01", "01", "00", "00", "11"),
262 => ("00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "01", "01"),
263 => ("01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "11", "11", "01", "01", "01"),
264 => ("00", "00", "11", "11", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "11", "01", "00", "00", "00"),
265 => ("00", "01", "00", "01", "01", "01", "11", "11", "00", "01", "00", "11", "01", "01", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01"),
266 => ("00", "00", "01", "00", "01", "11", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "11", "00", "01", "00"),
267 => ("01", "01", "01", "00", "11", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01"),
268 => ("00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "11", "11", "11", "01", "00", "00"),
269 => ("00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "11", "11", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01"),
270 => ("01", "00", "11", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00"),
271 => ("01", "00", "01", "11", "00", "00", "11", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "11", "00", "00", "01", "00"),
272 => ("00", "01", "11", "01", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00"),
273 => ("00", "00", "00", "11", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00"),
274 => ("01", "00", "01", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00"),
275 => ("01", "11", "00", "01", "00", "01", "01", "11", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01"),
276 => ("01", "00", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "11", "00", "11", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01"),
277 => ("01", "00", "01", "00", "00", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "01", "11", "00", "00", "01", "00", "11", "01", "00"),
278 => ("00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "11", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00"),
279 => ("00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "11", "00", "11", "01", "01", "11", "11", "00", "01"),
280 => ("00", "00", "00", "00", "00", "01", "01", "11", "00", "11", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "11", "00", "01"),
281 => ("01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "11", "00", "11", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "11", "01", "01", "01", "00"),
282 => ("01", "11", "00", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
283 => ("01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "11", "01", "11", "00", "11", "00", "00", "00", "00", "01", "01", "00"),
284 => ("01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "11", "00"),
285 => ("00", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "01", "11", "01", "00", "01", "01"),
286 => ("01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "11", "01", "11", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00"),
287 => ("00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "11", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00", "01", "11", "00", "00"),
288 => ("01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "11", "11", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11", "00", "00", "01", "01", "00"),
289 => ("00", "01", "11", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00"),
290 => ("01", "11", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01", "11", "00", "01", "01", "11", "01", "01"),
291 => ("00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "11", "11", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "11", "00", "01", "01", "00"),
292 => ("01", "01", "11", "01", "00", "01", "11", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01"),
293 => ("00", "01", "11", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "01"),
294 => ("01", "01", "00", "00", "00", "01", "11", "01", "01", "11", "00", "11", "11", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01"),
295 => ("00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "11", "01"),
296 => ("01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "11", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01"),
297 => ("01", "11", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "11", "01", "00", "01", "01", "11"),
298 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "11", "11", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "11", "00", "01"),
299 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "11", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11", "11"),
300 => ("00", "00", "11", "00", "01", "00", "01", "00", "11", "01", "11", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00"),
301 => ("01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "11", "00"),
302 => ("00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "11", "00", "11", "00", "01", "01", "01", "11", "11", "01", "00", "00", "00"),
303 => ("00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "11", "01", "00", "11", "01", "11", "01", "01", "00", "01", "01", "11"),
304 => ("00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "11", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "11"),
305 => ("00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "11", "01", "00", "11", "01", "00", "11", "01"),
306 => ("01", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00"),
307 => ("01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "11", "00", "01", "11", "00", "01", "01", "00", "00", "00"),
308 => ("01", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "01", "00", "11", "01", "11", "01", "00", "01", "01"),
309 => ("00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "01", "01", "00", "11", "01"),
310 => ("01", "11", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "11", "01", "11", "00", "01", "01", "01"),
311 => ("00", "00", "01", "11", "11", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "11", "01", "01", "11", "00", "00"),
312 => ("01", "01", "00", "01", "11", "01", "11", "00", "01", "11", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01"),
313 => ("01", "00", "11", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01"),
314 => ("00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "11", "01", "11", "00", "01"),
315 => ("01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "11", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "00", "11", "01", "00"),
316 => ("01", "01", "11", "01", "00", "11", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00"),
317 => ("01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "11", "01", "01"),
318 => ("01", "00", "01", "00", "11", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "01", "11", "00", "01", "01"),
319 => ("01", "00", "01", "11", "00", "00", "00", "00", "00", "11", "11", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01"),
320 => ("01", "00", "00", "11", "01", "00", "01", "00", "00", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00"),
321 => ("00", "11", "11", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01"),
322 => ("00", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "11", "01", "00", "00", "00"),
323 => ("00", "00", "11", "11", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "11", "11", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00"),
324 => ("00", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "11"),
325 => ("01", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00"),
326 => ("00", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "00", "11", "01", "11", "01"),
327 => ("01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11"),
328 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "11", "00", "01", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "11", "11", "01"),
329 => ("00", "00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00", "11", "00", "01", "00"),
330 => ("00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "00"),
331 => ("01", "00", "01", "11", "00", "01", "01", "01", "11", "11", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00"),
332 => ("01", "00", "01", "00", "00", "11", "01", "11", "01", "00", "00", "00", "01", "01", "11", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01"),
333 => ("00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "01"),
334 => ("00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "01", "11", "00", "01", "11", "01", "00", "11", "01", "01", "01", "00", "01"),
335 => ("00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "01", "11", "11", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01"),
336 => ("01", "01", "11", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00"),
337 => ("01", "00", "01", "00", "11", "11", "11", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
338 => ("00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "01", "00", "11", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00"),
339 => ("01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "01", "11", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "11", "01", "11"),
340 => ("01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "11", "11", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "11", "01", "00"),
341 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00"),
342 => ("01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "00", "11", "00", "00", "00", "11", "01", "00", "00"),
343 => ("00", "11", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01"),
344 => ("00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01", "11", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00"),
345 => ("01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "00", "11", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "11"),
346 => ("01", "11", "11", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00"),
347 => ("00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "11", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01"),
348 => ("01", "00", "01", "00", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11"),
349 => ("00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "11", "01", "01", "11", "01", "01", "01", "01", "00", "00", "11", "00"),
350 => ("01", "11", "00", "00", "11", "01", "00", "11", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00"),
351 => ("00", "01", "11", "00", "01", "01", "00", "11", "01", "00", "11", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00"),
352 => ("00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00"),
353 => ("00", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "00", "11", "01", "00", "00", "11", "00", "01", "01"),
354 => ("01", "01", "00", "00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "11", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01"),
355 => ("00", "01", "00", "01", "00", "00", "00", "11", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "11", "11", "01", "00", "00", "00", "01", "01", "00", "00"),
356 => ("01", "11", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00"),
357 => ("01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "00", "11", "00", "11", "00", "01", "00"),
358 => ("01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "11", "00", "11", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "00", "00"),
359 => ("01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "11", "00", "01", "11", "00", "11", "01", "01", "00"),
360 => ("01", "00", "11", "01", "00", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "11", "01", "00", "01", "01", "01", "01", "11"),
361 => ("01", "00", "00", "01", "00", "11", "11", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00"),
362 => ("01", "01", "00", "01", "01", "11", "01", "00", "11", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00"),
363 => ("01", "00", "01", "01", "00", "01", "01", "00", "11", "01", "11", "11", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01"),
364 => ("01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "11", "11", "01", "01", "11", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01"),
365 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "11"),
366 => ("00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "11", "01", "01", "01", "01"),
367 => ("01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11"),
368 => ("00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "11", "00", "00", "00", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "00"),
369 => ("01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "11", "00", "01", "01", "11", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "00"),
370 => ("01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01", "11", "00", "01", "00", "01", "01"),
371 => ("00", "11", "00", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "11", "11", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00"),
372 => ("00", "01", "11", "01", "00", "11", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "00", "00", "01"),
373 => ("01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "11", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01"),
374 => ("01", "01", "01", "11", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11", "01"),
375 => ("01", "00", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
376 => ("00", "01", "01", "00", "11", "00", "11", "01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00"),
377 => ("00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "11", "11", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01"),
378 => ("00", "01", "01", "01", "11", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "11", "00", "01", "01"),
379 => ("00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "11", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01"),
380 => ("01", "00", "00", "01", "11", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "01", "00", "11", "01", "01", "00", "00"),
381 => ("01", "00", "00", "01", "01", "11", "00", "11", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00"),
382 => ("00", "00", "01", "00", "00", "11", "01", "11", "11", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00"),
383 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "11", "00", "11"),
384 => ("00", "11", "01", "00", "11", "01", "11", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01"),
385 => ("01", "11", "00", "01", "00", "01", "01", "00", "11", "01", "11", "11", "11", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "01"),
386 => ("00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "11", "11", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00"),
387 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "11", "11", "00", "00"),
388 => ("01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "11", "11", "11", "00", "00", "00", "00", "01", "01"),
389 => ("00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "11", "00", "01", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "11", "00"),
390 => ("00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "11", "11", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00"),
391 => ("01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "11", "11", "01", "01", "11", "01", "01", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
392 => ("01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "00", "11", "00", "01", "00", "11", "01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "01"),
393 => ("00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "11", "00", "11", "01", "01", "11", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00"),
394 => ("01", "11", "01", "11", "00", "00", "00", "01", "01", "11", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01"),
395 => ("01", "00", "01", "11", "01", "00", "00", "11", "00", "00", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00"),
396 => ("01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01"),
397 => ("00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "11", "01", "11", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01"),
398 => ("00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "11", "01", "11", "00", "01", "00", "11", "01", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00"),
399 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "11", "11", "00", "00", "00", "00", "01", "00"),
400 => ("01", "01", "00", "01", "00", "01", "01", "11", "11", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "11", "11", "01", "01", "00", "00"),
401 => ("00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "11", "11", "11", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01"),
402 => ("01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "11", "01", "01", "00", "11", "11", "00", "00"),
403 => ("01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "11", "11", "00", "01", "01", "11", "01", "00"),
404 => ("01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "11", "01", "01", "11", "11", "00", "00", "01", "01"),
405 => ("01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "01", "11", "00", "00", "00", "11", "01", "00", "01", "00", "01", "01"),
406 => ("01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "11", "00", "01", "00", "01", "01", "00", "11", "11", "01", "00", "00", "00", "01", "00", "00"),
407 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "11", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "01", "11"),
408 => ("01", "11", "01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "11"),
409 => ("00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "11", "01", "11", "00", "01", "00", "00", "00", "01", "11", "11", "01", "00", "00", "00", "01", "01"),
410 => ("01", "01", "01", "00", "00", "00", "00", "11", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01"),
411 => ("00", "01", "00", "01", "01", "01", "11", "11", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "11", "00", "00", "00"),
412 => ("01", "01", "00", "01", "11", "01", "11", "00", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00"),
413 => ("00", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00"),
414 => ("00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "11", "01", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "11", "11"),
415 => ("01", "00", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00"),
416 => ("00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01"),
417 => ("00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "11", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00"),
418 => ("00", "01", "01", "01", "11", "00", "01", "11", "01", "11", "01", "00", "00", "01", "00", "00", "00", "11", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00"),
419 => ("00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "11", "01", "00", "11", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00"),
420 => ("01", "00", "01", "11", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "01", "01", "11", "01", "01", "00", "01", "11", "00"),
421 => ("00", "01", "11", "11", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01"),
422 => ("01", "11", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "01"),
423 => ("01", "11", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "00", "01", "11", "01", "01", "00", "01", "00", "01"),
424 => ("00", "11", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "11", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01"),
425 => ("00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "11", "11", "00"),
426 => ("01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "11", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11"),
427 => ("01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "11", "11", "01", "11", "00", "01", "00"),
428 => ("00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "11", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00"),
429 => ("00", "00", "11", "11", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00"),
430 => ("00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "11", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "11", "01", "11", "01", "01"),
431 => ("00", "11", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00"),
432 => ("01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "11", "01", "01", "01", "01", "01", "11", "01", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01"),
433 => ("00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "11", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01"),
434 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "11", "11", "00", "00", "00", "00", "01"),
435 => ("01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "00", "11"),
436 => ("00", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "11", "11", "01", "01"),
437 => ("01", "01", "00", "00", "11", "00", "01", "00", "01", "00", "11", "00", "01", "11", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01"),
438 => ("01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "11"),
439 => ("00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "11", "00", "11", "01", "01"),
440 => ("01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "11", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "11"),
441 => ("00", "00", "11", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01"),
442 => ("01", "00", "00", "01", "00", "01", "01", "01", "11", "11", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "11"),
443 => ("00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "11", "01", "11", "11", "01", "00", "01", "00", "01", "01", "01", "00"),
444 => ("00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "11", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
445 => ("01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "11", "01", "01", "01", "01", "00", "11", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01"),
446 => ("00", "00", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "00"),
447 => ("00", "00", "11", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00"),
448 => ("01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "00", "00", "11", "11", "01", "00", "01", "11", "00", "11", "01"),
449 => ("01", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "00", "11", "00", "00", "01", "01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
450 => ("00", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "11", "11", "00", "00", "01"),
451 => ("00", "00", "00", "00", "01", "01", "01", "00", "11", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "11", "01", "01", "01", "01"),
452 => ("00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "01", "11", "01", "11", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00"),
453 => ("00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "11", "01", "00", "11", "11", "00", "00", "01", "00", "11", "00"),
454 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "11", "01", "00", "01", "11", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "00"),
455 => ("01", "01", "00", "01", "00", "01", "00", "00", "11", "11", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01"),
456 => ("00", "01", "01", "11", "11", "00", "01", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01"),
457 => ("01", "00", "01", "00", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "00", "11", "01"),
458 => ("01", "00", "00", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00"),
459 => ("00", "01", "11", "01", "01", "01", "01", "00", "11", "11", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00"),
460 => ("01", "01", "01", "00", "00", "00", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01"),
461 => ("01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00"),
462 => ("01", "11", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00"),
463 => ("00", "01", "01", "11", "01", "11", "11", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00"),
464 => ("00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "11", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "11", "01"),
465 => ("00", "11", "11", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "00"),
466 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "11", "00", "11", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "11"),
467 => ("01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "11", "01", "11", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00"),
468 => ("01", "00", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "01", "11", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "11", "00", "01", "01"),
469 => ("00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "11", "01", "11", "00", "01", "11", "01", "01"),
470 => ("01", "11", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "11", "00", "11"),
471 => ("00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "11", "11", "01", "11", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00"),
472 => ("00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "00"),
473 => ("01", "00", "01", "11", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "11"),
474 => ("00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "00", "11", "11", "01", "01", "00"),
475 => ("01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "11"),
476 => ("01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "01", "00", "01", "00", "00", "11", "01"),
477 => ("01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "11", "01", "00", "01", "01", "11", "00", "11", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00"),
478 => ("00", "00", "00", "11", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "00"),
479 => ("00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "11", "00", "01", "00", "00"),
480 => ("00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "11", "11", "00", "11", "00", "00", "00"),
481 => ("00", "00", "00", "00", "01", "00", "11", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01"),
482 => ("00", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "00", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
483 => ("01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "11", "01"),
484 => ("01", "11", "01", "00", "11", "01", "11", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01"),
485 => ("01", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "11", "01", "00"),
486 => ("01", "01", "11", "11", "00", "11", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00"),
487 => ("00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "01", "11", "01", "01", "01"),
488 => ("00", "01", "11", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "01"),
489 => ("01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "11", "11", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
490 => ("01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01"),
491 => ("00", "00", "11", "11", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00"),
492 => ("01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "11", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01"),
493 => ("01", "01", "01", "01", "11", "00", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11"),
494 => ("00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "11", "00", "01", "00", "11", "00", "11"),
495 => ("01", "00", "11", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00"),
496 => ("01", "11", "00", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00"),
497 => ("01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "01", "11", "11", "00", "00"),
498 => ("01", "01", "01", "11", "00", "00", "00", "01", "01", "11", "00", "00", "11", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01"),
499 => ("01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "11", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "11", "01")),
(
0 => ("00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "11", "01", "11", "01", "01", "01", "01", "11", "01", "00"),
1 => ("00", "11", "11", "11", "00", "00", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "11", "00", "00", "00", "00"),
2 => ("01", "01", "00", "00", "01", "11", "00", "01", "00", "11", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00"),
3 => ("01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "11", "11", "01", "11", "00", "01", "11", "01"),
4 => ("00", "11", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11"),
5 => ("01", "01", "11", "01", "01", "11", "00", "00", "11", "01", "00", "00", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01"),
6 => ("00", "00", "01", "01", "00", "01", "01", "11", "11", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "11", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01"),
7 => ("00", "01", "00", "01", "00", "00", "00", "00", "11", "11", "11", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00"),
8 => ("00", "11", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "11", "00"),
9 => ("00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "11", "11", "11", "00", "11", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01"),
10 => ("01", "00", "00", "00", "01", "11", "01", "00", "11", "01", "00", "01", "11", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00"),
11 => ("01", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "11", "01", "11", "11", "01", "01", "00", "01", "00", "00", "01"),
12 => ("00", "00", "00", "11", "01", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "11", "11", "01"),
13 => ("01", "01", "01", "01", "11", "01", "01", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "11", "01"),
14 => ("00", "01", "00", "00", "11", "00", "00", "11", "01", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "01"),
15 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "11", "11", "00", "01", "01", "11", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00"),
16 => ("01", "00", "00", "01", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "11", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "11"),
17 => ("00", "00", "00", "00", "00", "01", "01", "01", "11", "11", "00", "01", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "11", "01", "01"),
18 => ("00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "11", "00", "11"),
19 => ("00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00", "11", "00", "01", "00", "01", "11", "00", "01", "11", "01", "01", "01", "00", "00", "11", "00", "00", "00", "11"),
20 => ("00", "01", "01", "11", "11", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00"),
21 => ("00", "01", "11", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "11", "00", "11", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00"),
22 => ("00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "11", "01", "00", "11", "01", "00", "01", "11", "11", "11", "01", "00", "00", "01"),
23 => ("00", "00", "00", "11", "00", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00"),
24 => ("01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "11", "11", "11", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01"),
25 => ("00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "11", "11", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "11"),
26 => ("01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "11", "11", "01", "11", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00"),
27 => ("01", "01", "01", "00", "00", "11", "00", "00", "11", "00", "11", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "11", "01", "11", "00", "01", "00", "00"),
28 => ("01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "11", "11", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01"),
29 => ("01", "01", "11", "01", "00", "01", "00", "11", "01", "11", "01", "00", "11", "00", "00", "01", "11", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "01"),
30 => ("01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "11", "01"),
31 => ("01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "11"),
32 => ("01", "11", "00", "11", "01", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "11", "01", "00", "00", "11", "00", "01", "00", "00", "00"),
33 => ("01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "11", "00", "11", "01", "01", "00", "11", "01", "00", "00"),
34 => ("00", "11", "00", "01", "01", "11", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "11", "01", "00", "11", "01", "01", "00", "00"),
35 => ("01", "00", "01", "11", "01", "00", "00", "00", "01", "11", "11", "00", "00", "11", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "01"),
36 => ("01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01", "00", "00", "00", "01", "11", "11", "01"),
37 => ("01", "01", "01", "01", "01", "01", "00", "11", "11", "11", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "11", "00"),
38 => ("01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01"),
39 => ("00", "11", "00", "00", "01", "11", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01"),
40 => ("01", "11", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "11", "00", "01", "00", "00", "00", "11", "01", "01", "11", "00", "00", "01", "01", "00"),
41 => ("00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "11", "01", "01", "01", "01", "11", "00", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00"),
42 => ("01", "00", "01", "11", "01", "00", "01", "11", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "01", "11", "01", "00", "11", "00"),
43 => ("00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "11", "00", "01", "00", "01", "01", "11", "00", "11", "00", "00", "00", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00"),
44 => ("01", "01", "01", "01", "11", "01", "11", "01", "01", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01"),
45 => ("01", "01", "00", "11", "01", "00", "11", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "00"),
46 => ("01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "11", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00"),
47 => ("01", "11", "01", "00", "00", "01", "11", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11"),
48 => ("00", "11", "01", "01", "01", "00", "01", "11", "00", "11", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01"),
49 => ("00", "00", "01", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00"),
50 => ("00", "11", "00", "01", "11", "11", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00"),
51 => ("00", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "11", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "11", "01", "11"),
52 => ("00", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "01", "00", "11", "01", "11", "11", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01"),
53 => ("01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "01", "00", "11", "01", "00", "11", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01"),
54 => ("00", "00", "01", "01", "11", "00", "00", "00", "01", "01", "11", "01", "11", "00", "01", "00", "11", "01", "00", "11", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00"),
55 => ("00", "11", "11", "00", "01", "11", "01", "11", "11", "01", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
56 => ("00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "11", "01", "11", "01", "00", "00", "01", "00", "11", "11", "00", "00"),
57 => ("00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "11", "11", "01", "00"),
58 => ("00", "01", "11", "00", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "00", "11"),
59 => ("00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "11", "01", "01", "00", "00"),
60 => ("01", "00", "11", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "11", "11", "01"),
61 => ("00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11", "01", "01", "11", "11", "01", "11", "00", "01", "01", "00", "00", "01", "11", "00", "00"),
62 => ("00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "01", "00", "11", "11", "01", "01", "11", "01", "01", "11", "00", "00"),
63 => ("00", "01", "11", "00", "01", "11", "11", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00"),
64 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "11", "00", "01", "00", "11", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "11"),
65 => ("01", "00", "00", "01", "00", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "11", "00", "00", "01", "00", "11", "01", "00", "00"),
66 => ("01", "00", "01", "11", "01", "01", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "11", "01", "01", "01", "11", "11", "00", "01", "01", "00", "01", "01", "01", "00", "01", "00"),
67 => ("00", "00", "01", "11", "00", "01", "11", "01", "11", "01", "00", "01", "00", "01", "00", "11", "00", "11", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
68 => ("00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "01", "11", "11", "00", "11", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01"),
69 => ("01", "11", "11", "11", "01", "00", "11", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
70 => ("01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "11", "00", "11", "00", "01", "01", "01", "01", "00", "11", "11", "01", "11", "00", "00", "00", "01"),
71 => ("01", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00", "11", "11", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
72 => ("00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "11", "11", "01", "01", "01", "11", "11", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01"),
73 => ("00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "00", "11", "00", "11", "01", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00"),
74 => ("01", "01", "01", "00", "00", "00", "01", "01", "00", "11", "11", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "11", "00", "00", "11", "00", "01"),
75 => ("00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "00", "11", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01"),
76 => ("00", "01", "01", "11", "00", "00", "00", "01", "11", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "01", "00", "11", "00"),
77 => ("00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01"),
78 => ("00", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "11", "01", "00", "00", "01", "11"),
79 => ("00", "11", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "11"),
80 => ("01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "11", "01", "00", "00", "11", "11", "01"),
81 => ("01", "01", "11", "11", "00", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
82 => ("00", "00", "00", "11", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "11"),
83 => ("00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "11", "00", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01"),
84 => ("00", "00", "11", "00", "11", "01", "00", "01", "00", "11", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01"),
85 => ("01", "01", "11", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "11", "11"),
86 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "01", "11", "11", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "11", "11", "01"),
87 => ("01", "11", "01", "11", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "11", "11", "00", "01"),
88 => ("00", "11", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "11", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00"),
89 => ("01", "00", "01", "00", "01", "11", "01", "01", "01", "11", "00", "11", "01", "01", "00", "11", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
90 => ("01", "00", "01", "11", "11", "01", "00", "00", "00", "00", "01", "01", "11", "11", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00"),
91 => ("00", "00", "00", "00", "01", "11", "01", "01", "01", "11", "01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00"),
92 => ("01", "01", "00", "01", "01", "01", "11", "11", "00", "00", "00", "11", "01", "11", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "01"),
93 => ("01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "11", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01"),
94 => ("00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "00", "00", "11", "01", "00", "00", "01", "11", "11"),
95 => ("01", "11", "00", "01", "00", "00", "11", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "01"),
96 => ("00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "11", "00", "01", "11", "01", "11", "00", "01", "11", "00", "00", "01", "00"),
97 => ("00", "11", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "11"),
98 => ("00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "00", "11"),
99 => ("00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "11", "11", "00", "00", "01", "00", "11", "11", "11", "01", "01", "01", "00", "00", "01"),
100 => ("01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "00", "11", "01", "11", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11"),
101 => ("01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "01", "01", "11", "00", "01", "11", "00", "00", "00", "00", "01", "00", "11", "01", "00"),
102 => ("00", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "11", "11", "00", "00"),
103 => ("01", "11", "11", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00"),
104 => ("01", "01", "11", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "01", "11", "01", "01", "00"),
105 => ("00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "11", "11", "00", "01", "11", "00", "00", "00"),
106 => ("00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "11", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "11", "01", "00"),
107 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "11", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "00", "11"),
108 => ("01", "11", "00", "01", "00", "01", "00", "11", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "11", "00", "01", "01", "01"),
109 => ("00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "11", "11", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11"),
110 => ("00", "01", "00", "00", "01", "00", "11", "11", "11", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00"),
111 => ("01", "00", "01", "00", "00", "11", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "11", "00"),
112 => ("00", "00", "11", "11", "00", "00", "00", "00", "01", "01", "11", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "01", "01", "00", "01", "00"),
113 => ("01", "11", "00", "00", "01", "11", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "11", "00"),
114 => ("01", "11", "01", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01"),
115 => ("00", "00", "00", "11", "00", "00", "01", "01", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00"),
116 => ("00", "11", "11", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11", "00"),
117 => ("00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "11", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00"),
118 => ("01", "11", "11", "11", "11", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00"),
119 => ("01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "11", "00", "01", "11", "00", "11", "00"),
120 => ("00", "00", "01", "11", "11", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "11"),
121 => ("01", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "11", "11", "01"),
122 => ("00", "11", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01"),
123 => ("01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "11", "01", "11", "01"),
124 => ("00", "11", "00", "00", "00", "00", "00", "11", "00", "01", "01", "11", "00", "11", "00", "00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01"),
125 => ("00", "01", "00", "11", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "01", "01", "11", "01", "11", "01"),
126 => ("01", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01", "11", "01", "01", "00", "11"),
127 => ("00", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "11", "01", "00", "00", "00", "01", "01", "11", "01", "11", "01"),
128 => ("01", "01", "00", "00", "01", "00", "11", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "11", "01", "11", "01", "00", "00", "11", "00", "00", "00", "01", "01"),
129 => ("00", "11", "11", "01", "00", "11", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00"),
130 => ("01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "00", "01", "00", "01", "11", "11", "00", "01", "00", "11", "01", "01", "11", "01", "01", "01", "11", "01", "01"),
131 => ("01", "01", "11", "00", "11", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "11", "01"),
132 => ("00", "11", "00", "01", "11", "11", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "11", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01"),
133 => ("00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "11", "00", "11", "01", "11", "00", "11", "01", "01", "01"),
134 => ("01", "00", "11", "11", "00", "01", "00", "11", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01"),
135 => ("00", "00", "01", "01", "00", "00", "11", "00", "00", "01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "11", "01", "00", "01", "01", "01", "11", "01", "00", "00"),
136 => ("01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "11", "00", "01", "00", "01", "00", "00"),
137 => ("01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "11", "01", "01", "11", "11", "01", "00", "11", "00"),
138 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11", "01", "01", "00", "00", "00", "00", "01", "11"),
139 => ("01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "11", "11", "01"),
140 => ("01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "11", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01"),
141 => ("01", "00", "01", "11", "01", "00", "01", "00", "01", "11", "01", "00", "11", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "00"),
142 => ("00", "00", "01", "01", "00", "11", "00", "01", "11", "00", "00", "01", "01", "11", "11", "11", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00"),
143 => ("00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "11"),
144 => ("00", "11", "01", "01", "00", "01", "00", "11", "11", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "11", "01", "01"),
145 => ("00", "01", "00", "11", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "11", "11", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01"),
146 => ("00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "11", "11", "00", "11", "01", "00", "01", "00", "01"),
147 => ("00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "00", "11", "00", "01", "01", "11", "00", "01", "00", "11", "00"),
148 => ("00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "11", "00", "01", "00", "11", "01", "01", "00", "11", "00", "01", "01"),
149 => ("01", "00", "00", "01", "11", "00", "01", "00", "00", "11", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "11"),
150 => ("00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01"),
151 => ("00", "11", "00", "01", "11", "00", "11", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "01"),
152 => ("01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "01", "00", "11", "01", "11", "01", "11", "00", "11", "01"),
153 => ("00", "00", "01", "00", "11", "00", "00", "11", "00", "01", "11", "01", "00", "01", "00", "11", "01", "11", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "00"),
154 => ("01", "01", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "11", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "11", "01", "00", "00"),
155 => ("00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "00", "00", "01", "11", "00", "11", "00", "00", "11", "11", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00"),
156 => ("01", "00", "11", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "11", "00", "01"),
157 => ("01", "01", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "11", "00", "00", "01", "00", "11", "00"),
158 => ("00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "11", "11", "01", "01", "00", "00", "01", "11", "01"),
159 => ("01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "01", "11", "11", "00", "00"),
160 => ("01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "11", "11", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11"),
161 => ("00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "01", "11", "00", "01", "01", "00", "01", "11", "00", "00", "11", "00", "00", "00", "11", "00", "00", "00", "11", "01"),
162 => ("01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "01", "00", "11", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11"),
163 => ("00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "01", "01", "00", "11", "01", "00", "00", "00", "11", "00", "00"),
164 => ("00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "11", "11", "01", "01", "01"),
165 => ("00", "00", "01", "11", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01", "11", "00", "01", "00", "00", "01", "00", "11", "00", "00", "01"),
166 => ("00", "11", "11", "00", "01", "01", "01", "01", "01", "11", "01", "11", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00"),
167 => ("00", "01", "11", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "11", "01"),
168 => ("00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "11", "11", "01", "00"),
169 => ("00", "01", "01", "11", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "11", "11", "01", "01", "00", "00", "00", "11", "01", "01", "01", "00"),
170 => ("00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "11", "01", "01", "11", "00", "00", "01", "11", "01", "11"),
171 => ("01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "11", "11", "01", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00"),
172 => ("00", "11", "01", "01", "11", "00", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "11", "01", "00", "01", "00", "00"),
173 => ("00", "01", "00", "11", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "00", "00", "00", "11", "11", "00", "00", "01", "01", "01", "00"),
174 => ("01", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "11", "00", "01", "01", "11", "00", "11", "11", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
175 => ("00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "00", "11", "01", "11", "01", "11", "00", "00", "00", "01", "00"),
176 => ("00", "11", "00", "11", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "11", "00", "00", "00"),
177 => ("00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "11", "11"),
178 => ("01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01"),
179 => ("01", "11", "01", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "11", "01", "00", "01", "11", "00", "00", "11", "00", "00", "01", "01"),
180 => ("01", "00", "00", "01", "11", "00", "11", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01", "11", "01", "01", "01", "00"),
181 => ("00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "11", "01", "01", "00", "11", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "00", "01"),
182 => ("00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "11", "00", "00", "00", "01", "00", "11", "01", "11", "01", "01", "00", "11"),
183 => ("01", "01", "11", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00"),
184 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "11", "00", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01", "11", "11", "00", "01", "11"),
185 => ("00", "01", "11", "00", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "01", "11"),
186 => ("01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "11", "01", "11", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "11", "01", "01", "00", "01"),
187 => ("00", "01", "00", "00", "00", "00", "11", "01", "11", "00", "00", "00", "00", "11", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00"),
188 => ("01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "11", "00", "01", "11", "01", "01", "11", "11", "01", "01", "01", "00", "00", "01", "00", "00"),
189 => ("01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "11", "11", "11", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "11"),
190 => ("00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "11", "00", "00", "00", "00", "11", "00", "01", "01", "11", "00", "11", "00", "00", "01"),
191 => ("01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "11", "00", "11", "01", "00", "00", "01", "00", "01", "11", "00"),
192 => ("01", "00", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "00", "11", "01", "11", "00", "00", "00", "00", "01", "01", "11", "00"),
193 => ("01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "11", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00"),
194 => ("00", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "11", "00", "11", "00", "00", "11", "11", "00", "00", "01", "00"),
195 => ("01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "11", "00", "00", "00", "00", "11", "00", "00", "11", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00"),
196 => ("00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11"),
197 => ("01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "01", "11", "00", "00", "11", "11", "00", "01", "01", "11", "00", "00"),
198 => ("01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00", "11", "00", "01", "11", "00", "01", "00", "01"),
199 => ("00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "11", "00", "00", "11", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01"),
200 => ("01", "00", "11", "00", "11", "11", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00"),
201 => ("00", "00", "11", "00", "01", "00", "01", "00", "11", "00", "11", "00", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "11", "01", "00"),
202 => ("01", "11", "00", "11", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "11", "01", "11", "00", "01", "00"),
203 => ("01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "11", "01", "00", "11", "01", "00", "00", "01", "11", "01"),
204 => ("01", "00", "01", "01", "11", "01", "01", "11", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00"),
205 => ("00", "01", "01", "00", "01", "00", "11", "01", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00", "11", "00", "00", "11", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
206 => ("00", "00", "01", "00", "11", "11", "00", "01", "00", "01", "00", "01", "11", "11", "00", "11", "00", "11", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00"),
207 => ("01", "11", "00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "11", "00", "11", "11", "01", "01", "00", "01"),
208 => ("01", "00", "01", "01", "00", "11", "11", "11", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00"),
209 => ("01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "11", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "01", "11", "00"),
210 => ("00", "11", "01", "01", "00", "00", "01", "00", "11", "11", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11"),
211 => ("00", "01", "01", "00", "00", "00", "00", "11", "11", "00", "01", "01", "11", "01", "01", "01", "11", "11", "11", "01", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00"),
212 => ("00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00", "11", "11", "01", "11", "01", "00"),
213 => ("00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "00", "11", "00", "00", "00", "00", "01", "00", "11", "11", "01", "00", "00", "01", "01", "01", "00", "11"),
214 => ("00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "11", "00", "11", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00"),
215 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "11", "01", "01", "11", "01", "00", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11"),
216 => ("00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "11"),
217 => ("00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "11", "00", "00", "11", "01", "00", "00"),
218 => ("01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "11", "00", "11", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00"),
219 => ("01", "01", "01", "00", "00", "01", "11", "11", "01", "11", "01", "01", "11", "01", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01"),
220 => ("00", "01", "01", "01", "01", "11", "00", "11", "01", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "11", "11", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01"),
221 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "01", "11", "11", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "11", "01", "00"),
222 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "11", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "00", "11", "00", "11", "01", "01", "01"),
223 => ("01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "11", "11", "01", "00", "00", "11", "01", "11", "01"),
224 => ("00", "00", "01", "11", "01", "00", "11", "01", "01", "01", "11", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00"),
225 => ("01", "11", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "11", "01", "01"),
226 => ("01", "11", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "01", "11", "00", "01", "11"),
227 => ("01", "01", "00", "00", "00", "01", "11", "01", "11", "01", "11", "01", "00", "01", "01", "11", "00", "00", "01", "00", "11", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01"),
228 => ("01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "01", "11", "00", "01", "00", "01", "11", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01"),
229 => ("01", "01", "11", "00", "01", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "11", "11", "00", "11", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01"),
230 => ("00", "01", "00", "11", "11", "00", "00", "11", "01", "11", "01", "01", "00", "00", "11", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00"),
231 => ("01", "00", "00", "00", "11", "00", "11", "00", "01", "00", "00", "11", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "11", "01", "01"),
232 => ("00", "01", "00", "01", "11", "00", "11", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "11", "00", "01", "00"),
233 => ("01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "11", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "11", "00", "11", "01", "00", "01", "01", "01", "01", "01"),
234 => ("00", "11", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "11", "11", "01", "01", "00", "00", "11", "01", "00", "01", "00", "00", "01", "11"),
235 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01"),
236 => ("01", "11", "01", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "11", "11", "00", "00", "01", "01", "00", "00", "01", "11", "00"),
237 => ("00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "00", "01", "11"),
238 => ("01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "00", "00", "11", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11"),
239 => ("00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "11", "00", "00", "11", "11", "01", "01", "00", "01", "11", "01", "01", "00", "11", "00", "01", "01", "00"),
240 => ("00", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "11", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00"),
241 => ("01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "01", "11", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11"),
242 => ("01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "11", "01", "11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "11", "01", "11", "01", "00", "00"),
243 => ("01", "00", "01", "11", "00", "00", "11", "01", "00", "01", "11", "01", "11", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "11"),
244 => ("00", "01", "11", "01", "01", "01", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "11", "11", "11", "01", "01"),
245 => ("01", "00", "01", "01", "00", "11", "00", "01", "11", "11", "01", "01", "00", "01", "11", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00"),
246 => ("00", "11", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "11", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01"),
247 => ("01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00", "11", "01", "11", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00"),
248 => ("00", "11", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "01", "00", "11", "01", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00", "01"),
249 => ("01", "01", "01", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "00", "11", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01"),
250 => ("00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "11", "00", "11"),
251 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "11", "01", "11", "11", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "01", "11", "01"),
252 => ("00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "11", "11", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "00", "11", "01"),
253 => ("01", "01", "00", "11", "01", "01", "00", "00", "01", "11", "11", "01", "00", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "11"),
254 => ("00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "00", "11", "00", "11", "01", "00", "00", "01", "11", "01", "11", "01", "00", "00"),
255 => ("00", "01", "11", "00", "00", "01", "11", "11", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01"),
256 => ("00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "11", "11", "00", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "11"),
257 => ("01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "11", "11", "11", "01", "11", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00"),
258 => ("00", "11", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01", "11", "00", "00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "00"),
259 => ("00", "00", "00", "00", "01", "01", "01", "00", "00", "11", "00", "11", "11", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "00"),
260 => ("01", "00", "01", "01", "11", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "00"),
261 => ("00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "11", "00"),
262 => ("00", "01", "11", "00", "00", "01", "11", "00", "01", "11", "01", "11", "01", "01", "11", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00"),
263 => ("01", "11", "11", "00", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "11", "01", "01", "01", "00"),
264 => ("00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "00", "11", "01", "11", "01", "01", "01", "00", "00", "11", "00", "01", "11", "00", "01", "00"),
265 => ("00", "11", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "01", "00", "11", "01"),
266 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "11", "00", "01", "00", "11", "00", "11", "01", "00", "01", "11", "00", "01", "01", "11", "01", "01"),
267 => ("01", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "11", "01", "11", "00", "01", "11", "11", "00", "00"),
268 => ("00", "01", "01", "00", "00", "00", "00", "11", "00", "11", "11", "00", "11", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01"),
269 => ("01", "00", "01", "01", "11", "11", "00", "11", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "11", "01", "01"),
270 => ("01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "11"),
271 => ("01", "01", "01", "00", "01", "01", "11", "11", "00", "01", "01", "11", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00"),
272 => ("00", "00", "01", "00", "00", "11", "00", "00", "01", "11", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "11", "01", "01", "11"),
273 => ("01", "01", "11", "00", "00", "01", "11", "00", "00", "00", "11", "00", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "11", "01"),
274 => ("01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "11", "00", "11", "00", "00", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00", "11", "01"),
275 => ("01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "11", "11", "01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00"),
276 => ("00", "01", "01", "11", "00", "01", "00", "01", "11", "11", "11", "00", "11", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "00"),
277 => ("01", "01", "01", "11", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00"),
278 => ("00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "11", "01", "11", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "01", "00", "00", "00"),
279 => ("00", "01", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "00", "00", "11", "01", "11", "01", "01", "11", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00"),
280 => ("01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "11", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00"),
281 => ("00", "01", "00", "11", "00", "00", "00", "01", "11", "00", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "11", "01", "00", "11", "00"),
282 => ("01", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "11", "01", "11", "01", "01", "01", "00", "01", "00"),
283 => ("00", "01", "01", "00", "01", "00", "00", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "11", "01", "01", "11", "01", "01"),
284 => ("01", "11", "00", "01", "11", "11", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "11", "00"),
285 => ("01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "11", "00", "01", "00", "00", "00", "11", "00", "01", "01", "11", "01", "00", "01", "00", "00", "11"),
286 => ("00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "11", "01", "11", "01", "11", "01", "11", "11", "01", "00"),
287 => ("01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "11", "00", "00", "00", "00"),
288 => ("01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "00", "01", "01", "00", "11", "11", "00", "01", "01", "01", "01", "01", "01", "00", "11", "11", "00", "00", "01", "01", "00", "00"),
289 => ("00", "01", "01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "01", "01", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00"),
290 => ("01", "00", "01", "11", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00"),
291 => ("00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "11", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "11", "01", "01", "01", "01", "01", "01"),
292 => ("01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "11", "01", "00", "00", "01", "11", "11", "00", "01", "01", "00", "00", "11", "11", "01", "01", "00"),
293 => ("01", "01", "00", "00", "01", "01", "11", "01", "11", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "11", "01", "11", "00", "00", "00", "01", "11", "01"),
294 => ("01", "01", "01", "01", "11", "01", "01", "11", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00"),
295 => ("00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "01", "11", "00", "01", "01", "01", "00", "01"),
296 => ("00", "00", "11", "00", "00", "11", "01", "01", "01", "00", "01", "01", "11", "01", "11", "01", "00", "01", "01", "11", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00"),
297 => ("01", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "11", "11", "01", "01", "01", "11", "00", "00", "11", "00", "01", "00", "01"),
298 => ("00", "01", "01", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "11", "01", "00"),
299 => ("01", "01", "00", "01", "11", "00", "01", "11", "11", "01", "11", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11"),
300 => ("01", "01", "11", "01", "01", "11", "11", "00", "01", "01", "11", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
301 => ("01", "01", "00", "01", "00", "11", "00", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00", "01", "11", "01", "11", "00", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
302 => ("01", "01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00", "01", "11", "00", "11", "11", "00", "01", "11", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01"),
303 => ("01", "11", "11", "01", "01", "00", "01", "11", "01", "11", "11", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00"),
304 => ("00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "11", "00", "11", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "11", "00", "00", "01", "11"),
305 => ("00", "00", "01", "01", "01", "01", "11", "11", "01", "11", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "11", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00"),
306 => ("01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "11", "00", "11", "00", "01", "11", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01"),
307 => ("01", "00", "11", "00", "11", "01", "00", "01", "11", "01", "11", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00"),
308 => ("01", "01", "00", "01", "01", "11", "01", "00", "11", "11", "11", "00", "11", "01", "00", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
309 => ("01", "11", "00", "01", "00", "00", "00", "11", "11", "00", "00", "11", "01", "11", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01"),
310 => ("00", "01", "00", "11", "11", "00", "01", "00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00"),
311 => ("00", "01", "11", "01", "11", "11", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00"),
312 => ("00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "11", "11", "01"),
313 => ("00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "01", "11", "01", "00", "01", "11", "01", "11", "00", "00", "00", "01", "01", "00", "00"),
314 => ("00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "11", "01", "01", "11", "11", "00"),
315 => ("00", "00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "11", "11", "00"),
316 => ("00", "00", "01", "00", "01", "01", "11", "01", "11", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "11"),
317 => ("00", "01", "01", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "11", "00", "11", "00", "01"),
318 => ("00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "11", "00", "00", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00"),
319 => ("00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "11", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "00", "01"),
320 => ("00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "11", "00", "11", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "11", "11", "00", "01"),
321 => ("00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "11", "11", "11", "01", "01", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "11", "00"),
322 => ("00", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "00", "11", "00", "00", "01", "00", "01", "11", "00", "01", "11", "11"),
323 => ("01", "00", "11", "00", "00", "01", "11", "01", "00", "01", "11", "11", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "01", "00", "00"),
324 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "11", "11", "00", "00", "01"),
325 => ("00", "11", "11", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11"),
326 => ("00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "11", "11", "01", "00", "00", "01", "00", "01", "00", "11", "11", "01", "00", "00", "01", "00", "01"),
327 => ("01", "11", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "11", "01", "01", "01", "11"),
328 => ("00", "00", "01", "11", "11", "00", "01", "00", "01", "11", "00", "11", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "01"),
329 => ("00", "01", "00", "11", "00", "00", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01"),
330 => ("00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "11", "01", "01", "00", "01", "00", "01", "11", "01", "11"),
331 => ("00", "11", "01", "00", "11", "01", "01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "01", "00", "11", "01"),
332 => ("00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "11", "00", "01", "11", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "11", "01"),
333 => ("00", "01", "01", "00", "01", "11", "00", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "11", "01", "00", "01", "00", "01", "01", "01"),
334 => ("01", "01", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00", "11", "01", "11", "11"),
335 => ("00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "00", "00", "00", "11", "00"),
336 => ("00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "11", "11", "00", "11", "00", "01", "00", "00", "11", "00", "01", "00"),
337 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "01", "11", "11", "01", "00"),
338 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "01", "00", "01", "11", "11", "11", "00", "00", "00", "01", "00", "11", "01", "00", "00"),
339 => ("01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "11", "00", "11", "01", "01", "11", "00", "01", "11", "01", "01", "01"),
340 => ("01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "11", "00", "11", "11", "01", "01", "01", "01"),
341 => ("00", "01", "00", "01", "00", "11", "00", "00", "00", "01", "11", "11", "00", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "11"),
342 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "11", "01", "01", "00", "00", "11", "11", "11", "01", "00", "01", "00", "00"),
343 => ("00", "01", "00", "11", "01", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "11", "01", "11", "01", "00", "01", "01"),
344 => ("00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "11", "01", "11", "01", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01"),
345 => ("00", "00", "01", "01", "00", "00", "11", "11", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "11", "00", "01"),
346 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "11", "01", "01", "01", "01", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
347 => ("01", "11", "01", "01", "11", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "00", "11", "01", "11", "01", "00", "01", "00"),
348 => ("00", "01", "00", "11", "11", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "11", "11", "01", "00", "01", "00", "01", "01", "00", "00"),
349 => ("00", "00", "01", "01", "00", "11", "00", "11", "01", "01", "00", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00"),
350 => ("01", "01", "11", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "01", "00", "01", "11", "11", "01", "01", "01", "00", "00", "00"),
351 => ("00", "01", "00", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "11", "00"),
352 => ("01", "00", "01", "11", "01", "00", "11", "11", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "01"),
353 => ("01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "11", "01", "11", "01"),
354 => ("01", "11", "00", "01", "11", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "11", "01", "11", "11", "00", "01", "00"),
355 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "00", "00", "11", "01", "01", "11", "01", "00"),
356 => ("01", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "11", "11", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "11", "00", "00", "00"),
357 => ("01", "01", "01", "11", "01", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "11", "11", "00"),
358 => ("00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "11", "01", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "11", "00", "01", "11", "01"),
359 => ("01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "01", "01", "11", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
360 => ("00", "01", "01", "11", "00", "01", "00", "00", "01", "11", "01", "01", "01", "00", "11", "11", "01", "00", "11", "00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00"),
361 => ("00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "11", "11", "00", "00", "01", "01", "00", "11", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "11", "01"),
362 => ("00", "00", "11", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "01"),
363 => ("01", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "00", "11", "00", "11", "11", "00", "00", "11", "00", "01", "01"),
364 => ("01", "11", "01", "00", "00", "01", "01", "11", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01"),
365 => ("01", "00", "00", "00", "01", "01", "11", "01", "00", "11", "11", "00", "11", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11"),
366 => ("01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "11", "00", "01", "01", "00", "11", "11", "00", "01", "11", "01", "11", "01", "00", "00", "00", "01"),
367 => ("00", "00", "00", "01", "00", "00", "01", "11", "11", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "01", "01"),
368 => ("00", "01", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "11", "01", "01", "11", "11", "11", "01", "01", "00", "00", "01"),
369 => ("01", "01", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "11", "11", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "00", "00"),
370 => ("01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "11", "01", "01", "01", "00", "01", "11", "00", "00", "11", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "11"),
371 => ("00", "11", "00", "01", "00", "00", "00", "11", "00", "00", "01", "11", "00", "01", "00", "00", "00", "11", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "11", "00", "00", "00"),
372 => ("00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "11", "01", "00", "01", "00", "01", "01", "11", "01", "01", "11", "01", "01", "11", "00", "01", "00", "00", "01", "00", "11"),
373 => ("01", "11", "11", "01", "11", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00"),
374 => ("00", "01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "11", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01"),
375 => ("00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "11", "00", "01", "11", "11", "00", "11", "00"),
376 => ("01", "00", "00", "00", "11", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "00", "00", "11", "01"),
377 => ("00", "11", "01", "00", "00", "11", "00", "01", "01", "11", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "11", "00", "00", "00", "01", "00", "00", "00"),
378 => ("01", "01", "00", "00", "01", "11", "11", "00", "00", "00", "01", "00", "01", "00", "00", "11", "11", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "01"),
379 => ("01", "11", "01", "01", "01", "00", "01", "11", "11", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01"),
380 => ("01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "11", "00", "00"),
381 => ("00", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "11", "00", "11", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01"),
382 => ("00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "11", "01", "01"),
383 => ("00", "01", "00", "01", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "01"),
384 => ("01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "11", "00", "01", "11", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "00", "11", "01", "01", "00", "11"),
385 => ("00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "11", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "11"),
386 => ("01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "11", "11", "00", "01", "01", "00", "01", "00", "11", "01", "11", "01"),
387 => ("00", "11", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01"),
388 => ("00", "00", "00", "11", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11"),
389 => ("00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "11", "11", "00", "01", "01", "01", "11", "01", "01", "11"),
390 => ("01", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "11", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "01", "11"),
391 => ("00", "11", "11", "00", "00", "01", "11", "00", "11", "00", "01", "01", "00", "11", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00"),
392 => ("01", "11", "11", "01", "00", "00", "01", "00", "11", "11", "00", "01", "01", "11", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
393 => ("00", "01", "01", "01", "01", "00", "11", "11", "01", "11", "00", "00", "00", "00", "01", "00", "11", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "01"),
394 => ("00", "11", "01", "00", "00", "00", "11", "01", "00", "11", "01", "11", "11", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01"),
395 => ("00", "11", "00", "00", "00", "11", "01", "01", "01", "00", "11", "01", "00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01"),
396 => ("00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "01", "00", "11", "11", "01", "00", "00", "01", "00", "11", "01", "01", "00", "00", "11", "01", "01", "01"),
397 => ("01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "11", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "11", "01", "01", "01", "01", "01", "11", "01", "01"),
398 => ("00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "11", "01", "11", "01", "01", "00", "01", "00", "11", "01"),
399 => ("01", "01", "11", "11", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "11"),
400 => ("01", "01", "00", "00", "00", "11", "00", "11", "01", "01", "01", "00", "01", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00"),
401 => ("01", "01", "00", "11", "00", "11", "11", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00"),
402 => ("00", "01", "01", "11", "00", "00", "11", "01", "01", "11", "01", "01", "01", "00", "00", "00", "01", "11", "11", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01"),
403 => ("00", "01", "01", "11", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "11", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00"),
404 => ("00", "01", "00", "01", "11", "11", "01", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00"),
405 => ("00", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "01", "00", "11", "00", "01", "01"),
406 => ("00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "11", "00", "00", "01", "01", "01", "11", "00", "11", "00"),
407 => ("00", "00", "00", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "01", "11", "00", "11", "01", "00", "11", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00"),
408 => ("01", "01", "11", "11", "11", "01", "11", "01", "00", "01", "00", "00", "01", "11", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00"),
409 => ("00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "11", "01", "00", "11", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "00", "11", "11"),
410 => ("00", "00", "11", "00", "01", "00", "11", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01"),
411 => ("01", "01", "01", "00", "01", "11", "00", "11", "00", "01", "11", "01", "00", "00", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11"),
412 => ("01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "00", "00", "00", "00"),
413 => ("00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "11", "00", "11", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01"),
414 => ("01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "11", "00", "00", "11", "00", "11", "00", "11", "01", "01", "01", "01", "01", "11", "01", "00"),
415 => ("00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "00", "01", "00", "01"),
416 => ("01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "00", "01", "11", "11", "01", "01", "00", "00", "11"),
417 => ("01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "11", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "01", "01", "00", "00", "00", "01", "00"),
418 => ("01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "11", "00", "00", "00", "00", "11", "01", "11", "00", "01", "01", "00", "00", "01"),
419 => ("01", "00", "01", "00", "00", "11", "00", "11", "11", "01", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "00", "01", "00"),
420 => ("01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "11", "11", "00", "11", "00", "01", "00", "00", "00", "01", "00"),
421 => ("00", "00", "01", "01", "01", "01", "11", "11", "01", "00", "00", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "11", "00"),
422 => ("00", "01", "00", "00", "00", "01", "11", "11", "01", "00", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01"),
423 => ("00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "11", "11", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "11", "00"),
424 => ("01", "00", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "11", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "11", "01", "00"),
425 => ("01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "01", "11", "01", "01", "11", "01", "00", "00", "00", "01", "11", "01", "01"),
426 => ("00", "11", "00", "11", "11", "00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
427 => ("01", "00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "01", "11", "00", "11", "11", "01", "01", "01", "01", "11", "00"),
428 => ("01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "11", "11", "00", "11", "00", "00", "00", "00"),
429 => ("01", "01", "00", "00", "00", "11", "11", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "11", "00", "01", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00"),
430 => ("01", "00", "01", "00", "01", "00", "00", "11", "01", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "11", "01", "11"),
431 => ("01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "11", "11", "01", "01", "11", "01", "01", "00"),
432 => ("01", "01", "01", "11", "11", "11", "11", "00", "01", "11", "00", "01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
433 => ("00", "01", "11", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "11", "11", "01", "01", "00", "00", "00", "11"),
434 => ("01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "01", "11", "01", "01", "11", "00", "00", "00", "00"),
435 => ("00", "00", "01", "01", "00", "00", "11", "11", "01", "11", "01", "11", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "00"),
436 => ("01", "01", "01", "01", "11", "01", "11", "11", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "00", "00", "01"),
437 => ("00", "00", "00", "01", "11", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "00", "11", "00", "00", "11", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "00"),
438 => ("00", "00", "11", "11", "01", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "01", "11", "11", "01", "01"),
439 => ("00", "00", "11", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11"),
440 => ("00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "11", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00"),
441 => ("01", "01", "01", "11", "01", "11", "00", "00", "00", "00", "11", "11", "00", "00", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00"),
442 => ("01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "11", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "11", "01"),
443 => ("01", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "00", "00", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "11", "01", "11"),
444 => ("00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "11", "11", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "00"),
445 => ("01", "01", "00", "11", "01", "11", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "01"),
446 => ("00", "00", "00", "00", "01", "11", "01", "00", "00", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "11", "11", "00", "01", "01", "00", "00", "01"),
447 => ("01", "01", "00", "01", "11", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "11", "11", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00"),
448 => ("01", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "11", "11", "11", "00", "01", "00", "00", "01"),
449 => ("01", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "00", "11", "00"),
450 => ("00", "01", "01", "01", "00", "01", "11", "00", "11", "01", "01", "01", "01", "11", "00", "01", "01", "00", "01", "11", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "00", "01"),
451 => ("00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "11", "01", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01"),
452 => ("00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00", "11"),
453 => ("01", "11", "01", "00", "00", "00", "00", "00", "00", "11", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00", "11", "00", "00"),
454 => ("01", "11", "01", "01", "01", "00", "11", "01", "00", "11", "00", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00"),
455 => ("01", "01", "00", "00", "01", "01", "11", "01", "01", "11", "00", "01", "01", "11", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "11"),
456 => ("00", "11", "11", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "11", "01", "11", "00", "01", "00", "01", "00", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
457 => ("00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "11", "01", "01", "00", "11", "00", "01", "00", "01", "11", "01", "11", "01", "01", "00", "00", "01", "01", "11", "01"),
458 => ("00", "11", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00"),
459 => ("01", "11", "00", "00", "01", "11", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "00"),
460 => ("01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "11"),
461 => ("00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "11", "01", "11", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00"),
462 => ("00", "11", "01", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "01", "01", "01", "01", "00", "11"),
463 => ("00", "00", "00", "11", "01", "01", "11", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00"),
464 => ("00", "00", "00", "01", "11", "01", "01", "01", "11", "01", "00", "11", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "11", "01", "01", "01", "00"),
465 => ("00", "11", "01", "00", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01"),
466 => ("01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "11", "11", "01", "01", "00", "01", "00", "00", "11", "01", "01", "11", "11", "01", "00"),
467 => ("01", "01", "01", "11", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "11", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01"),
468 => ("00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "11", "00", "11", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "11", "01"),
469 => ("01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "01", "11", "01", "11", "00", "00", "00", "00", "11", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00"),
470 => ("01", "00", "01", "11", "01", "00", "11", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "11"),
471 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11"),
472 => ("01", "00", "00", "00", "01", "01", "11", "00", "11", "11", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00"),
473 => ("01", "00", "00", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "11", "11", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01"),
474 => ("01", "11", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "00", "01", "11", "11", "00", "01", "01", "00", "01", "01"),
475 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00", "11", "00", "00", "11", "00", "00", "11", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00"),
476 => ("01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11", "00", "00", "00", "01"),
477 => ("01", "11", "01", "11", "00", "00", "00", "00", "01", "11", "00", "11", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00"),
478 => ("00", "01", "00", "00", "00", "11", "00", "01", "00", "11", "00", "01", "00", "11", "00", "11", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "00", "11", "00", "00", "01", "01"),
479 => ("01", "01", "01", "01", "11", "01", "11", "00", "01", "00", "01", "11", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "11", "01", "00", "01"),
480 => ("01", "00", "00", "01", "11", "00", "11", "01", "11", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00"),
481 => ("01", "11", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "01", "11", "00", "01", "11", "11", "01"),
482 => ("01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "11", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "00", "11", "00"),
483 => ("00", "00", "01", "11", "00", "01", "00", "01", "01", "11", "11", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "11", "01", "01", "01"),
484 => ("01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "11", "01", "01", "11", "00", "00", "01", "00", "11", "00"),
485 => ("00", "01", "00", "00", "11", "01", "00", "11", "11", "11", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00"),
486 => ("00", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00", "00", "11", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00"),
487 => ("01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "11", "11", "11"),
488 => ("00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "11"),
489 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "11", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "01", "01", "01"),
490 => ("01", "00", "00", "01", "00", "01", "11", "01", "00", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "11", "01", "00", "01"),
491 => ("01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "11", "01", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "00", "01", "00", "11", "11"),
492 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "11", "11", "00", "11", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "11"),
493 => ("01", "00", "01", "00", "00", "01", "01", "00", "11", "00", "00", "01", "11", "01", "11", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "11", "00", "00", "11", "01", "00", "00"),
494 => ("00", "00", "11", "00", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "00", "11", "01", "01", "00", "11", "00", "11", "00", "00", "00"),
495 => ("00", "11", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "01", "00", "01", "11", "01", "11", "11", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01"),
496 => ("01", "01", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "11", "00", "01", "11", "00", "11"),
497 => ("01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "11", "01", "01", "00", "01", "00", "01", "11", "11", "00", "00", "01", "11", "00", "11", "00", "00", "00"),
498 => ("01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "11", "11", "01", "00", "11", "11", "01", "01", "00"),
499 => ("01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "11", "11", "11", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00")),
(
0 => ("00", "01", "00", "11", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "11", "11", "01", "00", "01", "11", "01", "01", "00", "01"),
1 => ("00", "11", "01", "00", "11", "00", "01", "11", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "11", "00"),
2 => ("00", "01", "01", "00", "00", "11", "01", "00", "11", "01", "11", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "11", "00", "00"),
3 => ("00", "00", "01", "11", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00"),
4 => ("01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "11", "11", "01", "01", "11", "01", "00", "01", "00", "01", "01", "11"),
5 => ("00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "11", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "11"),
6 => ("01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "00", "00", "11", "01", "01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "11", "11", "00", "11", "01", "00", "00"),
7 => ("01", "01", "00", "11", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "01", "11", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01"),
8 => ("01", "11", "00", "01", "11", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "11"),
9 => ("00", "00", "00", "11", "00", "11", "00", "00", "01", "01", "01", "01", "11", "11", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "11", "00", "00", "11", "00", "01", "01"),
10 => ("01", "01", "00", "01", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "11", "11", "11", "00", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00"),
11 => ("01", "01", "11", "01", "11", "01", "00", "01", "11", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "00"),
12 => ("01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "11", "01", "11", "00", "01", "01", "11", "11", "01", "01", "11", "11", "00", "01", "01", "01", "00", "00", "01"),
13 => ("00", "01", "00", "00", "01", "11", "01", "11", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "11", "01", "00", "01", "11", "01", "11", "00"),
14 => ("00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01"),
15 => ("01", "01", "01", "01", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "11", "11", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "11", "00"),
16 => ("01", "01", "11", "11", "01", "00", "00", "00", "00", "00", "00", "11", "01", "11", "00", "01", "11", "01", "01", "00", "01", "11", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00"),
17 => ("01", "01", "01", "11", "01", "00", "11", "00", "01", "01", "11", "01", "11", "00", "00", "00", "00", "01", "00", "11", "00", "11", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01"),
18 => ("00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "11", "01", "01", "01", "00", "01", "01", "11", "00", "00", "00"),
19 => ("01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "11", "01", "00", "11", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "11", "01", "11"),
20 => ("00", "00", "11", "00", "01", "00", "00", "00", "11", "11", "11", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00"),
21 => ("00", "00", "00", "00", "11", "01", "11", "00", "01", "01", "11", "00", "00", "01", "00", "00", "01", "11", "11", "01", "11", "00", "01", "00", "01", "01", "01", "00", "01", "11", "00", "01"),
22 => ("00", "00", "11", "11", "11", "00", "01", "01", "01", "01", "00", "01", "11", "00", "11", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
23 => ("01", "01", "01", "11", "01", "11", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "11", "11"),
24 => ("00", "11", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "11", "00", "01", "01", "11", "11", "11"),
25 => ("00", "01", "00", "11", "11", "00", "01", "11", "00", "01", "11", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01"),
26 => ("01", "01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "01", "11", "11", "01", "00", "11", "11", "00", "11", "01", "11"),
27 => ("01", "01", "11", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "11", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "11", "01", "01", "00"),
28 => ("00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "00", "11", "00", "11", "00", "01"),
29 => ("00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "11", "11", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "11", "01", "00", "11", "01"),
30 => ("00", "01", "01", "00", "01", "01", "11", "11", "00", "11", "11", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "00", "11"),
31 => ("00", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "11", "11"),
32 => ("00", "00", "00", "00", "11", "11", "01", "00", "11", "01", "00", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "11", "01", "00", "11", "00", "01", "00", "11", "00", "00", "01"),
33 => ("01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "11", "11", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "11", "00", "01", "01", "11", "01", "11"),
34 => ("01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "11", "01", "01", "01", "01", "11", "00", "01", "00", "11", "01", "11", "00", "01", "01", "00", "11", "01"),
35 => ("01", "01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "00", "11", "01", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "11"),
36 => ("01", "00", "01", "11", "11", "11", "00", "11", "00", "11", "11", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01"),
37 => ("01", "01", "01", "00", "01", "11", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "00", "11", "00", "01", "01", "00", "11", "00", "11", "00", "00"),
38 => ("01", "01", "00", "01", "11", "00", "01", "01", "01", "00", "11", "01", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "11", "00", "00", "11", "01", "00", "11", "11", "00", "01"),
39 => ("01", "11", "01", "00", "00", "00", "00", "01", "00", "11", "01", "11", "01", "11", "11", "00", "00", "00", "00", "01", "11", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "01"),
40 => ("01", "11", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "11", "11", "00"),
41 => ("01", "00", "11", "01", "00", "11", "11", "01", "00", "00", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "11", "01", "01", "01", "00"),
42 => ("01", "01", "00", "01", "01", "00", "00", "11", "11", "01", "00", "00", "11", "01", "00", "00", "11", "00", "01", "01", "11", "01", "00", "11", "00", "11", "00", "00", "00", "00", "01", "00"),
43 => ("01", "01", "01", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "11", "01", "11", "00", "00", "11", "11", "01", "01", "11", "11", "00", "00", "01", "00", "00", "00"),
44 => ("00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "11", "00", "00", "11", "11", "01", "01", "11", "11", "00", "00", "00", "01", "01", "01", "00", "11"),
45 => ("01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "11", "11", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "11"),
46 => ("01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "00", "11", "11", "00", "01", "00"),
47 => ("00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "11", "00", "11", "11", "01", "11", "00", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "01"),
48 => ("01", "11", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "11"),
49 => ("00", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "00", "11", "11", "00", "01", "01", "11", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00"),
50 => ("01", "01", "11", "11", "01", "00", "11", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "00", "01"),
51 => ("01", "01", "11", "01", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "11", "01", "00", "11", "01"),
52 => ("00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "11", "11", "11", "00", "00", "01", "00", "01", "01", "00", "01", "11"),
53 => ("01", "01", "11", "00", "01", "00", "00", "11", "01", "00", "01", "01", "11", "01", "11", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11"),
54 => ("00", "00", "11", "00", "00", "00", "11", "11", "11", "00", "00", "00", "11", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "00"),
55 => ("00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "11", "00", "01", "11", "01", "11", "01", "01", "00", "00", "11", "01", "01"),
56 => ("00", "11", "00", "01", "01", "00", "01", "01", "00", "00", "11", "11", "11", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "00", "01", "00"),
57 => ("01", "11", "00", "00", "11", "01", "11", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "11", "01", "00", "00", "00", "00", "11", "11", "00", "00", "01", "00", "01", "01"),
58 => ("01", "11", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "11", "01"),
59 => ("01", "01", "01", "11", "01", "11", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "11"),
60 => ("00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "01", "11", "11", "00", "11", "01", "01"),
61 => ("01", "01", "00", "00", "00", "00", "01", "11", "01", "01", "11", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "11"),
62 => ("00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "01", "11", "01", "11", "01", "11", "01", "01", "11", "01", "00"),
63 => ("00", "11", "11", "11", "11", "01", "01", "01", "00", "11", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11"),
64 => ("01", "01", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "11", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01"),
65 => ("00", "11", "11", "00", "01", "11", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "11", "11", "01", "01", "01", "11", "00"),
66 => ("01", "01", "01", "01", "01", "01", "11", "11", "01", "00", "11", "01", "00", "01", "01", "00", "11", "11", "01", "01", "11", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "01"),
67 => ("01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "11", "00", "00", "01", "00", "01", "11", "00", "01", "01", "11", "00", "11", "00", "11", "01", "11", "00", "01", "00", "01", "01"),
68 => ("00", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "00", "11", "11", "00", "01", "11", "01"),
69 => ("00", "11", "01", "01", "00", "01", "11", "01", "00", "11", "01", "00", "11", "00", "01", "00", "00", "11", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11"),
70 => ("00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "11", "01", "00", "01", "11", "00", "01", "00"),
71 => ("01", "00", "00", "01", "00", "11", "00", "01", "11", "01", "01", "11", "01", "00", "01", "11", "00", "00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "00"),
72 => ("00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "00", "01", "11", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "11", "00", "01", "00", "01", "00"),
73 => ("01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "01", "11", "01", "01", "11", "01", "11", "01", "00", "11", "00", "01", "01", "11", "01", "00", "01", "01"),
74 => ("01", "00", "01", "11", "00", "01", "11", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "11", "11", "00", "01", "00", "00", "11", "00"),
75 => ("01", "00", "01", "01", "01", "01", "11", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "11", "01", "00", "01", "11", "00", "01", "11", "01", "01", "00", "01"),
76 => ("01", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "11", "11", "01", "01", "00", "11", "00", "01", "01", "11", "00", "11", "01", "01", "01"),
77 => ("00", "01", "00", "00", "11", "00", "01", "00", "01", "11", "00", "11", "01", "00", "00", "11", "00", "00", "11", "00", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01", "11", "01"),
78 => ("00", "00", "00", "01", "11", "00", "11", "01", "11", "00", "00", "01", "00", "11", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01"),
79 => ("01", "11", "01", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "11", "00", "00", "11", "01", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01"),
80 => ("00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "11", "00", "11", "01", "11", "11", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "11", "01", "01", "00"),
81 => ("00", "00", "01", "11", "11", "11", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "11", "00", "01", "11", "00", "00"),
82 => ("00", "11", "00", "01", "00", "11", "01", "00", "11", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01"),
83 => ("01", "01", "00", "11", "01", "00", "01", "11", "00", "01", "00", "11", "01", "01", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "11", "00", "00", "11", "00"),
84 => ("01", "00", "00", "11", "11", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01"),
85 => ("01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "00", "01", "11", "00", "01", "00", "00"),
86 => ("00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "11", "11", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "01", "00"),
87 => ("00", "01", "01", "11", "11", "11", "01", "11", "01", "11", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00"),
88 => ("01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "11", "00", "00", "11", "00", "00", "00", "11", "01", "11", "00", "11", "01", "01", "00", "00"),
89 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "01", "11", "11", "00", "00", "00", "00", "11", "11", "00", "01", "11", "01", "11", "01", "01", "01"),
90 => ("00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "11", "01", "00", "11", "11", "01", "00", "11", "00", "01", "01"),
91 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "11", "11", "11", "01", "01", "01", "11", "01", "01", "00"),
92 => ("00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "01", "11", "00", "00", "00", "11", "11", "01", "11", "11", "01", "01", "00", "01"),
93 => ("01", "01", "00", "11", "01", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "11", "00", "00", "00", "11", "00"),
94 => ("00", "11", "11", "00", "11", "11", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01"),
95 => ("01", "00", "01", "00", "11", "00", "00", "00", "00", "00", "11", "00", "11", "01", "01", "11", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "11", "11", "00"),
96 => ("00", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "11", "11", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11"),
97 => ("01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "11", "01", "11", "00", "01", "11", "00", "01", "00"),
98 => ("00", "00", "01", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "11", "01", "11", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11", "01", "00", "11", "00", "01"),
99 => ("00", "01", "01", "01", "01", "01", "11", "11", "00", "00", "01", "01", "00", "01", "00", "11", "11", "11", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "00"),
100 => ("00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "01", "01", "11", "01", "01", "00", "11", "01", "01", "01", "11", "01", "00", "00", "11", "01", "11", "00", "11", "01"),
101 => ("00", "01", "11", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "11", "01", "11", "01", "00", "00", "01", "11", "00", "01"),
102 => ("00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "00", "00", "11", "00", "00", "11"),
103 => ("00", "01", "00", "11", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "00", "11", "01"),
104 => ("00", "00", "01", "11", "00", "00", "11", "01", "01", "11", "00", "11", "01", "11", "01", "00", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11"),
105 => ("01", "00", "01", "11", "00", "01", "01", "11", "01", "00", "00", "00", "11", "01", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "11", "01", "01", "01"),
106 => ("00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "00", "00", "11", "11", "00", "00", "01", "11", "01", "01", "11", "01"),
107 => ("01", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01"),
108 => ("00", "00", "01", "01", "01", "00", "11", "00", "00", "11", "00", "01", "01", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "11", "00"),
109 => ("01", "00", "11", "11", "00", "00", "11", "01", "00", "00", "11", "01", "00", "00", "00", "00", "01", "11", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01"),
110 => ("01", "01", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "11", "01", "01", "00", "01", "00", "11", "00", "11", "11", "00", "01", "11", "01", "00", "00", "01", "01"),
111 => ("00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "11", "01", "11", "11", "01", "01", "00", "11", "11", "01", "01", "01", "00", "01"),
112 => ("01", "00", "00", "01", "01", "11", "01", "00", "00", "11", "11", "00", "01", "00", "01", "01", "01", "11", "00", "11", "01", "01", "11", "11", "00", "01", "01", "00", "00", "00", "00", "01"),
113 => ("00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "11"),
114 => ("00", "01", "11", "01", "00", "01", "00", "01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "11", "01", "01", "11", "00", "00", "11", "00"),
115 => ("00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "01", "11", "01", "11", "01", "00", "00", "11", "00", "00", "11", "00", "00", "01", "01", "01"),
116 => ("00", "00", "01", "00", "00", "00", "11", "01", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "01", "11", "00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01"),
117 => ("00", "00", "01", "11", "01", "01", "11", "01", "00", "00", "11", "01", "00", "11", "01", "01", "00", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11"),
118 => ("00", "01", "00", "00", "11", "01", "11", "00", "00", "00", "11", "11", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "11", "00", "11"),
119 => ("00", "00", "11", "01", "01", "11", "01", "11", "11", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00"),
120 => ("01", "01", "01", "01", "01", "01", "00", "01", "11", "00", "11", "01", "11", "01", "01", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00"),
121 => ("01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "11", "00", "00", "01", "11", "01", "11"),
122 => ("01", "01", "01", "00", "01", "00", "01", "01", "11", "11", "11", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "11", "00", "11"),
123 => ("01", "01", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "11", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "11"),
124 => ("01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "00", "11", "01", "01", "00", "01", "11", "11", "00", "01", "01", "01", "00", "11", "00", "01", "00", "11", "01", "01", "11"),
125 => ("00", "01", "00", "00", "00", "01", "01", "11", "01", "00", "11", "00", "01", "11", "00", "01", "01", "00", "00", "01", "11", "01", "01", "11", "01", "00", "11", "01", "01", "00", "01", "00"),
126 => ("00", "11", "00", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "00", "01", "01", "00", "11", "01", "11"),
127 => ("01", "01", "01", "11", "11", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "11", "01", "00", "01", "00", "01", "01", "11", "11", "00", "01"),
128 => ("00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "11", "11", "11", "01", "01", "11", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00"),
129 => ("00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "11", "01", "11", "11", "01", "01", "01", "00", "01", "00", "00", "11"),
130 => ("01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "01", "01", "11", "11", "00", "01"),
131 => ("01", "01", "01", "11", "11", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "11", "01", "00", "00", "01", "11", "00", "11", "01"),
132 => ("01", "01", "01", "00", "01", "00", "00", "01", "11", "11", "01", "11", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01"),
133 => ("00", "01", "11", "01", "00", "11", "00", "11", "11", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "00"),
134 => ("01", "01", "00", "11", "00", "11", "00", "00", "00", "00", "00", "01", "11", "01", "11", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00"),
135 => ("00", "00", "00", "01", "00", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "11", "01", "01", "01", "01", "00", "00", "11", "11", "00", "00", "11", "01"),
136 => ("01", "01", "01", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "11", "11", "11", "11", "01", "01", "00", "00", "00", "01"),
137 => ("00", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "11", "11", "00", "11", "01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "11"),
138 => ("00", "11", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "11", "11", "01", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01"),
139 => ("01", "01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "00", "11", "11", "00", "11", "01", "00", "00", "11"),
140 => ("00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "11", "01", "11", "00", "01", "01", "00", "11", "00", "01", "11", "01"),
141 => ("01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "01", "11", "01", "00", "11", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "11", "11", "01", "01", "00"),
142 => ("01", "11", "01", "00", "00", "00", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "11", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "11", "00", "00"),
143 => ("00", "11", "00", "11", "00", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "11", "11", "01", "01", "00", "00"),
144 => ("00", "00", "00", "00", "01", "11", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "01", "01", "01"),
145 => ("01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "01", "11", "11", "00", "00", "01", "11", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "11", "11", "01"),
146 => ("00", "11", "11", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "11", "01", "01", "01", "01", "11", "00"),
147 => ("01", "00", "11", "01", "01", "01", "11", "01", "00", "11", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00", "00", "01", "11", "01", "01", "00"),
148 => ("00", "00", "00", "01", "01", "11", "11", "00", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "11", "01"),
149 => ("00", "11", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "11", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00"),
150 => ("00", "11", "11", "11", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00"),
151 => ("01", "00", "11", "00", "00", "01", "01", "01", "11", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "11", "00", "11", "01", "01", "01", "00", "11", "01", "01"),
152 => ("00", "11", "11", "00", "00", "00", "01", "00", "00", "01", "11", "00", "00", "00", "11", "01", "00", "11", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "01"),
153 => ("01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "01", "11", "11", "11", "01", "11", "00", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "11", "01", "01", "00"),
154 => ("01", "00", "00", "01", "00", "00", "01", "11", "00", "00", "11", "00", "01", "00", "00", "01", "11", "00", "11", "01", "01", "00", "01", "00", "11", "00", "00", "00", "11", "00", "01", "11"),
155 => ("01", "00", "01", "01", "00", "00", "11", "01", "11", "01", "11", "00", "01", "01", "11", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00"),
156 => ("01", "11", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "00", "11", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00"),
157 => ("00", "11", "11", "01", "01", "01", "11", "01", "00", "01", "00", "11", "11", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "11", "00", "01", "00", "00", "00", "00"),
158 => ("00", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "11", "11", "00", "11", "01", "00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "00", "00", "01", "00"),
159 => ("01", "00", "00", "00", "00", "01", "00", "11", "11", "00", "01", "00", "11", "01", "11", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "00", "11"),
160 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "11", "11", "01", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "01", "00", "11", "00", "01"),
161 => ("01", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "01", "01", "11", "00", "11", "00", "00", "11", "11", "01", "01", "11", "01", "01", "11", "00"),
162 => ("00", "00", "01", "11", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "11", "01", "01", "01", "11"),
163 => ("00", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "00", "11", "00", "11", "01", "01", "11", "01", "01", "00", "11", "01", "00", "01"),
164 => ("01", "01", "01", "00", "01", "11", "11", "01", "00", "00", "00", "11", "11", "11", "01", "00", "11", "01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00"),
165 => ("00", "00", "00", "11", "01", "11", "01", "11", "01", "00", "00", "01", "00", "01", "11", "11", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "01", "01", "00", "01", "00", "00"),
166 => ("01", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "11", "11", "00", "11", "00", "11", "01", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00"),
167 => ("00", "00", "00", "11", "00", "01", "11", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "11", "00", "11", "01", "11", "01", "11", "00", "00", "00"),
168 => ("01", "01", "01", "00", "00", "00", "11", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "11", "01", "01", "11", "00", "00", "11", "00", "01", "11"),
169 => ("01", "01", "00", "11", "11", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "11", "00", "11", "01", "11", "01", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01"),
170 => ("00", "11", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "11"),
171 => ("00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "11", "00", "01", "11", "00", "11", "01", "00", "00", "00", "01", "11", "00", "01", "00", "01"),
172 => ("00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "11", "00", "00", "01", "11", "01", "11", "01", "00"),
173 => ("00", "00", "00", "00", "01", "11", "11", "11", "00", "11", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "11", "01"),
174 => ("00", "00", "01", "11", "00", "01", "00", "11", "01", "11", "01", "00", "01", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00", "11"),
175 => ("00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "11", "11", "11", "01", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "11", "00", "01", "11"),
176 => ("00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "11", "11", "01", "00", "00", "01", "11", "01", "01", "11", "01", "11", "00", "00", "00", "00", "00", "01", "01"),
177 => ("00", "00", "01", "00", "00", "00", "11", "01", "11", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "11", "11", "00", "00", "00", "01"),
178 => ("00", "00", "11", "01", "11", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01"),
179 => ("01", "11", "00", "01", "00", "11", "01", "00", "00", "00", "00", "00", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "11", "11", "01", "00", "01", "01", "01", "11"),
180 => ("01", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "11", "01", "00", "11", "01", "01", "00", "11", "11", "01", "01", "00", "00", "11", "01", "00", "11", "00", "00"),
181 => ("01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "11", "11", "11", "00", "11", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01"),
182 => ("00", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00", "00", "11", "11", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01"),
183 => ("00", "11", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "11", "11", "11", "01", "01", "00"),
184 => ("00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "11", "11", "00", "11", "00", "01", "01", "11"),
185 => ("00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "11", "11", "00", "00", "00", "01", "11", "01", "11", "00", "00"),
186 => ("00", "00", "00", "11", "01", "00", "00", "01", "01", "11", "00", "00", "11", "01", "00", "00", "01", "00", "11", "00", "01", "11", "00", "11", "01", "01", "01", "11", "01", "00", "00", "00"),
187 => ("01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "00", "11", "00", "00", "01", "11", "01"),
188 => ("00", "00", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "11", "11", "00", "11", "00", "01", "00"),
189 => ("01", "00", "01", "01", "01", "01", "11", "00", "11", "00", "01", "01", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "11", "11", "01"),
190 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "11", "11", "01", "11", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00"),
191 => ("01", "11", "00", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "11", "01"),
192 => ("00", "00", "00", "11", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "11", "01", "00", "00", "11", "01", "11", "00", "11", "00"),
193 => ("01", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "11", "00", "00", "11", "11", "11", "11"),
194 => ("00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "11", "01", "01", "11", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "11"),
195 => ("01", "00", "01", "01", "00", "11", "00", "00", "01", "11", "00", "11", "01", "11", "11", "00", "01", "00", "01", "01", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00"),
196 => ("00", "00", "11", "00", "00", "11", "00", "01", "00", "11", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "00", "11", "00", "11"),
197 => ("00", "00", "00", "01", "11", "00", "11", "00", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "00"),
198 => ("01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "11", "11", "11", "11", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
199 => ("00", "00", "00", "01", "01", "01", "11", "11", "00", "11", "01", "00", "01", "01", "01", "01", "11", "00", "00", "11", "01", "00", "00", "11", "01", "01", "01", "00", "01", "00", "11", "01"),
200 => ("01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "11", "11", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "11", "11"),
201 => ("01", "01", "11", "00", "00", "00", "01", "11", "11", "11", "01", "01", "11", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "00"),
202 => ("01", "00", "11", "00", "11", "01", "11", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "01", "00", "11"),
203 => ("01", "01", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "11", "11", "01", "11", "01", "01", "11", "01", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "00"),
204 => ("01", "01", "00", "01", "01", "00", "01", "11", "01", "11", "01", "00", "11", "00", "00", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "11", "00", "11", "01", "01", "11"),
205 => ("00", "11", "11", "00", "00", "11", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00"),
206 => ("01", "11", "00", "01", "00", "11", "11", "00", "01", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "11", "00", "11", "00", "00"),
207 => ("00", "11", "00", "00", "11", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "00"),
208 => ("00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "11", "01", "11", "00", "11", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01"),
209 => ("01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "11", "11", "00", "11", "11", "01", "01", "01", "01", "00", "01", "11", "00"),
210 => ("01", "00", "11", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "11", "01", "00", "00", "01", "01", "01", "00", "11", "11", "01", "01", "00", "11"),
211 => ("01", "01", "00", "11", "01", "11", "00", "11", "11", "01", "01", "01", "01", "01", "11", "11", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "00"),
212 => ("01", "00", "00", "01", "11", "00", "00", "00", "11", "11", "11", "11", "01", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00"),
213 => ("00", "00", "00", "00", "01", "00", "00", "11", "01", "11", "01", "11", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11", "01", "11", "01", "01", "01"),
214 => ("00", "01", "01", "00", "11", "01", "11", "00", "01", "00", "01", "01", "11", "11", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "01", "00", "11", "11", "00"),
215 => ("01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "00", "00", "11", "11", "01", "01", "11", "01"),
216 => ("00", "00", "01", "01", "00", "01", "11", "11", "01", "11", "00", "00", "11", "00", "11", "00", "00", "11", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "01", "01", "01"),
217 => ("01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "11", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "00", "11", "01", "11", "00", "01", "11"),
218 => ("00", "11", "11", "00", "00", "11", "00", "11", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00"),
219 => ("00", "11", "01", "11", "00", "00", "11", "01", "01", "00", "11", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00"),
220 => ("01", "11", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "11", "11", "00", "00"),
221 => ("01", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "11", "11", "00", "01"),
222 => ("00", "00", "00", "00", "00", "00", "00", "11", "11", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "11", "01", "01", "01", "11", "01", "01", "11", "00", "00", "11", "00", "01"),
223 => ("01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "11", "11", "00", "00", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "11", "01", "01", "01"),
224 => ("01", "11", "00", "01", "00", "01", "11", "01", "00", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00"),
225 => ("00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "11", "11", "11", "00", "01", "01", "00", "01", "01", "11", "11", "00", "01", "00", "00", "00", "11"),
226 => ("01", "00", "00", "11", "11", "00", "00", "11", "00", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "00", "11", "00", "11", "00", "01", "01", "01", "00", "01", "11", "00"),
227 => ("01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "00", "11", "11", "01", "11", "01", "01", "00", "00", "11", "01", "00", "00", "01", "11", "11", "00", "00", "01", "00", "00"),
228 => ("00", "01", "01", "11", "00", "11", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00"),
229 => ("01", "00", "01", "11", "00", "01", "01", "00", "01", "11", "00", "00", "11", "11", "00", "11", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00"),
230 => ("00", "01", "00", "00", "11", "11", "11", "11", "11", "01", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01"),
231 => ("00", "01", "01", "00", "11", "00", "11", "11", "01", "11", "11", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "11", "01", "01", "01", "01", "01"),
232 => ("00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "00", "11", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "01", "11", "11", "11"),
233 => ("01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "11", "01", "11", "01", "01", "00", "11", "00", "11", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01"),
234 => ("00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "00", "11", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "11", "01", "00", "11", "00", "11"),
235 => ("01", "00", "01", "01", "00", "11", "00", "00", "11", "00", "00", "11", "01", "01", "11", "01", "01", "01", "01", "00", "11", "11", "01", "01", "11", "01", "00", "00", "01", "00", "01", "01"),
236 => ("00", "00", "01", "00", "11", "01", "00", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "11", "01", "01", "11", "01", "00", "00", "01", "01", "11", "01", "11"),
237 => ("01", "00", "11", "11", "00", "00", "00", "01", "11", "00", "01", "11", "11", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01"),
238 => ("01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "11", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "11", "11", "11", "11", "01", "01", "01", "01", "01"),
239 => ("00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "11", "11", "01", "00", "11", "11", "01", "01", "00", "01", "01", "00", "11"),
240 => ("01", "11", "11", "11", "11", "01", "00", "01", "11", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00"),
241 => ("01", "00", "00", "01", "00", "01", "00", "11", "11", "01", "11", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "11", "01", "00", "11", "00", "01"),
242 => ("01", "11", "01", "11", "11", "01", "01", "01", "01", "01", "11", "00", "11", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01"),
243 => ("00", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "00", "11", "01", "00", "11", "11", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "01"),
244 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "11", "11", "00", "01", "01", "11", "01", "00", "11", "11", "00", "11", "00", "01", "01", "01", "01", "01", "00", "01"),
245 => ("00", "01", "00", "01", "00", "11", "01", "00", "11", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "01", "11", "01", "01"),
246 => ("00", "01", "00", "11", "00", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "00", "01", "01", "00", "11", "00", "11", "00", "11", "00", "00", "11", "00", "01", "01", "00", "01"),
247 => ("00", "00", "01", "01", "11", "00", "00", "11", "11", "00", "00", "01", "00", "00", "11", "01", "00", "11", "11", "01", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "01"),
248 => ("00", "11", "11", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00"),
249 => ("01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "11", "11", "01", "00", "11"),
250 => ("00", "00", "01", "00", "00", "00", "01", "11", "01", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "11", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00"),
251 => ("01", "01", "01", "01", "00", "11", "01", "11", "01", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "11", "01", "01", "11", "11"),
252 => ("00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "11", "11", "00", "11", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "11", "01"),
253 => ("00", "00", "01", "01", "01", "00", "11", "00", "00", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "00", "11", "01", "00", "11", "11", "00", "00"),
254 => ("01", "11", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "11", "00", "00", "00", "11", "00", "11", "00", "01"),
255 => ("01", "00", "11", "01", "00", "01", "01", "11", "01", "01", "01", "01", "11", "11", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "00"),
256 => ("00", "01", "11", "11", "00", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "11", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "01", "01"),
257 => ("01", "11", "11", "11", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "11", "00", "00", "00", "00"),
258 => ("00", "01", "00", "11", "00", "01", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "11", "01", "01"),
259 => ("00", "01", "00", "01", "11", "00", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "01", "11", "11", "01"),
260 => ("01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "11", "11", "11", "01", "01", "01", "01", "00", "11"),
261 => ("01", "01", "11", "00", "01", "01", "00", "00", "11", "11", "00", "01", "01", "11", "00", "01", "01", "00", "01", "01", "11", "11", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00"),
262 => ("01", "11", "01", "00", "00", "11", "01", "11", "00", "11", "01", "00", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00"),
263 => ("00", "01", "01", "11", "01", "01", "11", "00", "00", "00", "01", "01", "01", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "11", "00", "01", "00", "01"),
264 => ("01", "11", "00", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "11", "01", "11", "01", "01", "01"),
265 => ("00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "11", "11", "00", "00", "01", "00", "00", "11", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11"),
266 => ("01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "00", "01", "11"),
267 => ("01", "01", "00", "11", "00", "00", "11", "00", "01", "11", "11", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "00", "01", "11", "00", "01", "00"),
268 => ("01", "01", "01", "00", "11", "11", "11", "00", "01", "00", "00", "01", "00", "00", "11", "00", "11", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01"),
269 => ("00", "00", "00", "01", "01", "01", "11", "00", "01", "01", "11", "00", "11", "11", "00", "00", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "00", "01", "01", "01"),
270 => ("01", "01", "11", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "01", "01", "11", "01", "00", "01", "01", "01", "11", "01", "00", "11", "01", "11"),
271 => ("01", "01", "00", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "00", "00", "00"),
272 => ("01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "01", "01", "11", "00", "01", "11", "11", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00"),
273 => ("00", "01", "01", "00", "11", "11", "01", "01", "01", "11", "01", "01", "01", "01", "11", "01", "11", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01"),
274 => ("01", "00", "01", "01", "00", "11", "00", "01", "11", "00", "01", "01", "01", "00", "01", "11", "00", "01", "00", "01", "11", "01", "01", "01", "01", "01", "01", "00", "01", "11", "11", "00"),
275 => ("00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "11", "00", "11", "01", "01", "11", "01", "01", "11"),
276 => ("01", "00", "01", "11", "01", "01", "01", "11", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "01", "11", "00", "01", "11", "11", "01"),
277 => ("00", "00", "00", "11", "00", "01", "01", "01", "01", "11", "11", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "11", "01", "01", "11"),
278 => ("01", "00", "00", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "11", "01", "01", "01", "11", "11", "00", "11"),
279 => ("00", "11", "00", "11", "00", "00", "01", "11", "00", "01", "01", "11", "00", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00"),
280 => ("01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "11", "00", "01", "01", "11", "00", "00", "00", "01", "00", "11", "00", "11", "00", "00", "01", "01"),
281 => ("01", "11", "00", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "11", "00", "11", "11", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "01"),
282 => ("00", "00", "00", "00", "01", "01", "11", "01", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "11", "11", "00", "11", "01", "01", "00"),
283 => ("01", "01", "00", "00", "01", "11", "01", "00", "01", "01", "11", "00", "00", "00", "11", "01", "11", "01", "00", "01", "11", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00"),
284 => ("01", "00", "11", "01", "11", "00", "11", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01", "11"),
285 => ("01", "00", "11", "11", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "00", "11", "11", "01", "11", "01", "01", "00", "00", "00", "00", "01"),
286 => ("00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "01", "01", "11", "11", "11", "01", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "11", "00", "11", "01", "01"),
287 => ("01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "11", "00", "00", "01", "00", "11", "11", "11", "00", "11", "01", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01"),
288 => ("01", "00", "01", "11", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "11", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "01", "11"),
289 => ("01", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "11", "11", "11", "01", "11", "01", "01", "00", "00", "01", "01", "11", "01"),
290 => ("00", "11", "01", "11", "01", "01", "01", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01"),
291 => ("00", "00", "01", "00", "11", "00", "11", "01", "01", "11", "01", "11", "11", "11", "01", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "01"),
292 => ("01", "11", "00", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01", "11", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01"),
293 => ("00", "11", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "01", "00", "11", "01", "00", "01", "11", "00", "11", "01"),
294 => ("01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00", "11", "00", "00", "01", "11"),
295 => ("01", "01", "00", "01", "00", "11", "11", "01", "01", "11", "01", "00", "00", "11", "00", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "00", "11", "01", "01", "01"),
296 => ("01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "11", "00", "01", "00", "01", "01", "11", "01", "11", "01", "00", "01", "11", "00", "00", "01", "11"),
297 => ("01", "00", "00", "01", "01", "01", "11", "01", "11", "00", "00", "11", "11", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11"),
298 => ("01", "01", "01", "11", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00"),
299 => ("01", "00", "00", "11", "01", "00", "00", "00", "00", "11", "00", "00", "11", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "00"),
300 => ("00", "01", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "11", "01", "11", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00"),
301 => ("00", "11", "01", "00", "01", "11", "00", "00", "00", "00", "01", "11", "00", "00", "01", "00", "01", "00", "11", "11", "01", "11", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00"),
302 => ("01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "00"),
303 => ("00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "11", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "00", "01", "11", "00", "00"),
304 => ("00", "01", "11", "01", "00", "00", "00", "01", "11", "01", "01", "11", "01", "00", "11", "11", "01", "00", "00", "01", "11", "01", "00", "11", "01", "00", "00", "01", "01", "00", "01", "00"),
305 => ("01", "11", "11", "00", "11", "01", "01", "01", "00", "11", "11", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "01"),
306 => ("01", "00", "01", "11", "01", "01", "11", "11", "00", "00", "01", "11", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "11", "00", "00"),
307 => ("01", "00", "00", "01", "11", "01", "00", "01", "11", "01", "01", "00", "11", "01", "11", "00", "11", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "00", "01", "00"),
308 => ("01", "00", "00", "01", "01", "00", "11", "01", "11", "01", "11", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00", "00", "11"),
309 => ("00", "01", "01", "00", "00", "11", "01", "11", "11", "01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "00", "01", "00"),
310 => ("01", "01", "01", "00", "11", "01", "01", "01", "01", "00", "00", "11", "11", "11", "01", "00", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "11", "01"),
311 => ("01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "11", "01", "00", "11", "01", "01", "11", "01", "01", "00", "00", "01", "11", "01", "00", "01", "11", "00", "01", "01", "01", "01"),
312 => ("01", "01", "00", "00", "00", "00", "11", "00", "11", "00", "01", "11", "00", "00", "00", "11", "01", "11", "00", "01", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "00"),
313 => ("00", "11", "00", "00", "00", "11", "00", "00", "01", "11", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "00", "11", "01", "11", "01", "00"),
314 => ("01", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "00", "11", "01", "00", "11", "00", "00", "01", "00", "00", "00", "11", "11", "11", "01", "00", "00", "00", "01", "01", "01"),
315 => ("00", "00", "00", "11", "01", "00", "11", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11", "00"),
316 => ("01", "00", "00", "00", "00", "11", "01", "11", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "00", "11", "11", "00", "01"),
317 => ("00", "11", "01", "11", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "00", "11", "00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00"),
318 => ("00", "11", "00", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "11", "00", "01", "11", "00", "01", "00", "00", "11", "00", "01", "01", "11", "01", "01", "01", "01", "11"),
319 => ("01", "01", "00", "11", "11", "11", "00", "11", "01", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00"),
320 => ("01", "11", "00", "11", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "11", "11", "11", "00", "00", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00"),
321 => ("00", "11", "00", "00", "11", "00", "00", "11", "11", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "01", "01", "01", "01", "00", "11", "00", "00", "00", "01"),
322 => ("00", "01", "00", "01", "11", "00", "01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "11", "11", "01", "01", "01", "01", "01", "01"),
323 => ("00", "01", "00", "00", "00", "00", "01", "11", "11", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "01", "11", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01"),
324 => ("01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "11", "00", "01", "11", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01"),
325 => ("01", "01", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "00", "11", "00", "00", "11", "01", "11", "00", "11", "00", "00", "01", "00", "11"),
326 => ("00", "11", "01", "00", "00", "00", "01", "11", "01", "00", "11", "11", "01", "01", "00", "00", "01", "01", "01", "00", "01", "00", "11", "11", "00", "00", "11", "01", "00", "01", "00", "00"),
327 => ("00", "01", "00", "00", "11", "00", "00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "11", "00", "00", "00", "01", "11", "11", "00", "00", "11", "01", "00", "01", "01", "00"),
328 => ("00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "00", "00", "01", "00", "11", "11", "00", "00"),
329 => ("00", "00", "01", "01", "11", "11", "01", "01", "01", "11", "11", "01", "00", "01", "00", "11", "00", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "01"),
330 => ("01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "00", "01", "01", "00", "11", "00", "11", "00", "00", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "11", "00", "11"),
331 => ("00", "01", "00", "00", "00", "11", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11"),
332 => ("00", "11", "01", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01", "11", "11", "11", "01", "01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00"),
333 => ("00", "00", "01", "11", "01", "00", "00", "00", "11", "00", "00", "11", "11", "00", "01", "00", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00"),
334 => ("00", "00", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "01", "11"),
335 => ("00", "00", "01", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "11", "00", "11", "11", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "00"),
336 => ("01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "00", "11", "11", "00", "01", "11", "01", "11", "01", "01"),
337 => ("00", "00", "11", "01", "00", "01", "01", "11", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "11", "01", "01", "01", "11", "01", "00", "01"),
338 => ("00", "01", "01", "11", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "11", "01", "01", "11", "00"),
339 => ("01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "11", "11", "01", "00", "01", "00", "11", "11", "00", "01", "00", "01", "00"),
340 => ("00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "11", "01", "11", "01", "01", "11", "01", "01"),
341 => ("00", "00", "00", "01", "01", "11", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "11", "11", "00", "01", "11", "11", "01", "01", "11"),
342 => ("00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "11", "01", "11", "00", "01", "01", "01", "01", "00", "01", "11", "11", "11", "01", "01", "00", "01", "01", "00"),
343 => ("00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "01", "11", "01", "11", "11", "00", "11", "00", "01"),
344 => ("00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "11", "11", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "11", "00", "00", "11", "01"),
345 => ("00", "00", "11", "11", "11", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "11", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "01", "01"),
346 => ("01", "11", "01", "00", "01", "01", "00", "11", "11", "11", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01"),
347 => ("00", "11", "01", "11", "01", "00", "01", "11", "00", "01", "00", "11", "01", "01", "11", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01"),
348 => ("01", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "11", "11", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "11", "11", "00", "00"),
349 => ("01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "11", "00", "01", "01", "11", "11", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "01"),
350 => ("01", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "01", "01", "00", "11", "01", "01", "11", "11", "00", "11", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01"),
351 => ("00", "11", "00", "11", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "00", "11", "01", "11", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "11"),
352 => ("00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "01", "11", "11", "01", "00", "00", "11", "11", "01", "01", "01", "00", "01", "11", "00", "00", "11", "01", "01", "01"),
353 => ("01", "01", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "01", "11", "11", "11", "00", "01", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01"),
354 => ("00", "00", "01", "01", "00", "11", "11", "00", "01", "01", "11", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "00", "11", "11", "00", "00", "00", "11", "00", "00", "00"),
355 => ("01", "01", "01", "11", "01", "11", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00"),
356 => ("01", "01", "01", "00", "00", "11", "00", "11", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "11", "11", "11", "00", "00"),
357 => ("00", "01", "01", "11", "00", "01", "01", "01", "01", "11", "01", "01", "00", "11", "11", "01", "11", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "11", "01"),
358 => ("01", "01", "00", "00", "00", "11", "00", "01", "11", "00", "01", "01", "00", "01", "01", "01", "11", "01", "11", "00", "11", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "00"),
359 => ("01", "00", "01", "11", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "01"),
360 => ("00", "11", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "11", "00", "11", "00", "01", "11", "11", "00", "00", "00", "00", "01", "00", "01"),
361 => ("00", "01", "11", "00", "00", "01", "11", "01", "01", "00", "01", "11", "01", "11", "00", "11", "11", "00", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "01"),
362 => ("01", "11", "11", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "11", "00", "11"),
363 => ("00", "00", "11", "00", "00", "11", "01", "01", "01", "01", "00", "00", "11", "11", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01"),
364 => ("00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "11"),
365 => ("00", "11", "11", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01", "11", "11", "00", "00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "11", "01", "00", "00"),
366 => ("00", "00", "01", "01", "00", "01", "00", "01", "01", "11", "11", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "11", "00", "00", "01", "01"),
367 => ("00", "01", "01", "00", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "11", "00", "11", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01"),
368 => ("00", "01", "11", "00", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "11", "01", "00", "11", "00", "11", "00", "01", "01", "00", "00", "01", "00"),
369 => ("01", "01", "11", "00", "11", "11", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01"),
370 => ("00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "01", "11", "11", "00", "11", "00", "00", "01"),
371 => ("01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "00", "11", "11", "01", "00", "00", "11", "00", "01"),
372 => ("01", "00", "01", "01", "00", "11", "01", "11", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "00", "11", "11", "01", "11", "00", "11", "00", "01", "00", "00", "01", "01"),
373 => ("00", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00", "01", "11", "01", "01", "11", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "11"),
374 => ("00", "01", "00", "11", "01", "01", "01", "11", "01", "00", "01", "01", "01", "00", "11", "11", "11", "00", "01", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "01", "11"),
375 => ("00", "01", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "11", "01", "01", "11", "00", "00", "00", "01", "01", "11"),
376 => ("00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "11", "11", "00", "00", "01", "00", "01", "00", "00"),
377 => ("01", "11", "01", "11", "11", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "11", "11", "00", "01", "01"),
378 => ("00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "11", "01", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "00", "11", "11", "01", "00", "11", "01", "01"),
379 => ("01", "00", "11", "01", "00", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "11", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "01", "00"),
380 => ("01", "01", "11", "01", "01", "11", "11", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "11", "00"),
381 => ("00", "00", "11", "11", "01", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "11", "11", "01", "00", "01", "11", "00", "01", "01", "01", "00", "01"),
382 => ("01", "00", "11", "11", "00", "01", "00", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "11", "11", "00", "00", "01"),
383 => ("01", "00", "01", "00", "11", "01", "00", "01", "11", "00", "00", "11", "01", "01", "00", "11", "01", "00", "01", "01", "00", "00", "01", "01", "01", "11", "00", "11", "01", "01", "00", "11"),
384 => ("01", "11", "01", "00", "11", "00", "00", "00", "01", "11", "11", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01"),
385 => ("00", "00", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "11", "01", "01", "00", "00", "11", "11", "11", "00", "00", "00"),
386 => ("00", "01", "11", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "11", "00", "11", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "11", "00"),
387 => ("01", "00", "01", "11", "01", "00", "11", "11", "00", "01", "00", "00", "00", "00", "01", "00", "11", "11", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "01", "01"),
388 => ("01", "00", "01", "11", "11", "00", "01", "11", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "11", "00", "01", "00", "01"),
389 => ("00", "01", "01", "11", "11", "00", "11", "11", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "00"),
390 => ("01", "00", "01", "11", "00", "01", "01", "11", "01", "11", "11", "01", "00", "00", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "00", "00", "00", "01"),
391 => ("00", "11", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "11", "00", "00", "11", "11", "00", "00", "01", "11", "01"),
392 => ("01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "01", "00", "01", "01", "01", "00", "11", "11", "01", "00", "01", "01", "00", "11", "00", "11", "00", "00", "00"),
393 => ("01", "00", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "11", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "11", "00", "00", "01", "00", "11"),
394 => ("00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00", "11", "00", "11", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "11", "01", "00"),
395 => ("01", "00", "01", "11", "11", "01", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "01", "11", "01", "01", "01", "01", "00", "11", "01", "01", "01", "11", "00"),
396 => ("00", "00", "00", "11", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "01", "11", "11", "11", "00", "11", "00", "00", "11", "00", "00", "00", "00"),
397 => ("00", "01", "00", "01", "01", "00", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "11", "01"),
398 => ("01", "11", "00", "01", "01", "01", "11", "00", "11", "00", "00", "00", "01", "01", "00", "11", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00"),
399 => ("01", "11", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "11", "00", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00"),
400 => ("00", "01", "00", "11", "01", "11", "00", "00", "11", "00", "00", "01", "01", "11", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00"),
401 => ("00", "01", "00", "01", "11", "01", "01", "11", "00", "11", "00", "00", "01", "11", "01", "00", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "11", "01", "01", "11"),
402 => ("00", "01", "01", "00", "01", "00", "11", "00", "01", "01", "01", "11", "00", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "01", "11", "11"),
403 => ("01", "00", "01", "00", "11", "00", "00", "01", "00", "01", "11", "11", "11", "00", "11", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "11", "00"),
404 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "11", "00", "01", "00", "00", "11", "01", "00", "01", "00", "11", "01", "11", "11"),
405 => ("01", "01", "01", "01", "00", "00", "11", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "11", "00", "11", "11", "01", "11", "00", "01"),
406 => ("01", "01", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "00", "11", "01", "11", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "11"),
407 => ("01", "01", "00", "01", "11", "11", "00", "00", "01", "00", "11", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "01"),
408 => ("00", "00", "11", "11", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00"),
409 => ("01", "01", "01", "11", "00", "01", "01", "11", "11", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "01", "01", "01", "00", "11"),
410 => ("01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01", "00", "11", "00", "01", "11", "01"),
411 => ("00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "11", "11", "01", "01", "11", "01", "00", "00", "01", "11", "00", "01", "01"),
412 => ("01", "11", "00", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "11", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00"),
413 => ("01", "00", "01", "01", "00", "11", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "01", "01", "01", "00", "11", "00", "01", "01", "11", "00", "11", "00", "01", "11"),
414 => ("00", "01", "00", "00", "11", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11"),
415 => ("01", "00", "00", "00", "00", "11", "01", "01", "11", "01", "00", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "11", "00", "00", "00", "00", "11", "01", "00"),
416 => ("01", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "11", "11", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00"),
417 => ("00", "01", "01", "01", "11", "00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "11", "00", "00", "01", "01", "11", "01", "01", "00", "11", "11"),
418 => ("00", "11", "00", "00", "11", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "11", "01", "11", "00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00"),
419 => ("00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "00", "11", "00", "01", "00", "11", "00", "01", "11", "00", "01", "00"),
420 => ("00", "00", "11", "00", "00", "11", "00", "01", "01", "00", "11", "01", "00", "01", "00", "11", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00"),
421 => ("00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "00", "11", "11", "11", "11", "01", "01", "00"),
422 => ("00", "01", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "11", "01", "11", "01", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11", "11", "00", "11", "00", "01"),
423 => ("00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "11", "00", "01", "00", "11", "01", "01", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01"),
424 => ("00", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "11", "11", "11", "00", "00", "11", "00", "01", "00", "01", "00", "11", "01", "00", "00", "00"),
425 => ("00", "00", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "00", "01", "01", "11", "11", "01", "00", "11", "01", "11", "00", "00", "11", "00", "11", "01", "00"),
426 => ("00", "01", "00", "01", "11", "01", "01", "00", "11", "11", "00", "11", "01", "01", "01", "01", "01", "01", "01", "01", "00", "11", "11", "01", "11", "00", "01", "00", "01", "00", "01", "01"),
427 => ("00", "11", "01", "00", "00", "01", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "11", "00", "01", "11", "01", "01"),
428 => ("00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01", "11", "00", "00", "00", "11", "01", "11", "01", "00", "11", "01", "00", "11", "01"),
429 => ("01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "11", "00", "11", "00", "01", "01", "11", "01", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "11", "00", "01"),
430 => ("00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "00", "11", "01", "00", "11", "01", "01", "01", "11", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "00", "00"),
431 => ("01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "00", "11", "00", "00", "01", "01", "01", "00", "11", "00", "11", "11", "00", "00", "01", "01", "00"),
432 => ("00", "01", "11", "01", "11", "01", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "11"),
433 => ("01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00", "01", "00", "01", "00", "00", "11", "11", "11", "00", "11", "11", "00", "00", "00", "00"),
434 => ("00", "01", "11", "00", "01", "01", "11", "01", "01", "01", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "11", "11", "00", "00", "11", "01"),
435 => ("01", "11", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "11", "11", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01"),
436 => ("01", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "01", "01", "00", "11", "11", "11", "01", "00", "11", "01", "11", "11", "01", "01"),
437 => ("01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "11", "11", "00", "01", "00", "01", "01", "00", "11"),
438 => ("00", "01", "00", "01", "00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "11", "00", "01", "11", "01", "00", "01", "01", "00", "01", "11", "00", "11", "00", "11", "01", "11"),
439 => ("00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "11", "11", "01", "11", "01", "00", "11", "00", "11", "01", "01", "01"),
440 => ("00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "11", "11", "11", "01", "00", "11", "01", "01", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01"),
441 => ("00", "11", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "00", "11", "00"),
442 => ("01", "11", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "01", "11", "11", "00", "11", "00"),
443 => ("00", "01", "00", "11", "11", "00", "00", "01", "11", "00", "00", "00", "00", "00", "11", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "01"),
444 => ("01", "01", "01", "01", "01", "11", "01", "01", "00", "11", "11", "01", "01", "00", "11", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "00"),
445 => ("00", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "11", "01", "00", "11", "00", "00", "11", "00", "00", "01", "00", "11", "01"),
446 => ("00", "01", "01", "01", "11", "11", "01", "00", "01", "11", "00", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00"),
447 => ("00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "11", "11", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
448 => ("01", "11", "00", "11", "01", "11", "00", "11", "11", "01", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "00"),
449 => ("01", "00", "00", "00", "00", "11", "11", "11", "00", "01", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "11"),
450 => ("00", "11", "01", "01", "01", "00", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "00", "01", "00", "01", "11", "00"),
451 => ("00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11", "01", "11", "01", "11", "00", "00", "00", "11", "11", "01", "01", "01", "00", "00", "00", "01", "01"),
452 => ("00", "11", "00", "01", "01", "01", "11", "01", "00", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "11", "11", "01"),
453 => ("00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "11", "00", "01", "11", "11", "00", "01", "01", "01", "01", "00", "00", "00", "11", "11", "01", "01", "01", "00", "01", "00", "01"),
454 => ("01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11", "11", "00", "00", "00", "11"),
455 => ("01", "01", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "00", "00", "11", "11", "00", "00", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "11"),
456 => ("00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "11", "01", "11", "11", "00", "01", "11", "00", "01", "01", "01", "11", "00"),
457 => ("00", "11", "11", "00", "00", "11", "00", "01", "00", "11", "00", "00", "11", "01", "01", "01", "11", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "01"),
458 => ("00", "01", "11", "11", "00", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "11", "01", "01", "11", "01", "00", "01", "01", "01"),
459 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "11", "00", "00", "00", "11", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00", "01", "11"),
460 => ("01", "11", "00", "00", "01", "01", "00", "11", "00", "00", "11", "11", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00", "11"),
461 => ("01", "01", "01", "00", "01", "01", "01", "11", "11", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "11", "01", "11", "01", "00", "01", "00", "01", "00", "11"),
462 => ("01", "11", "01", "11", "00", "01", "01", "00", "01", "00", "00", "11", "00", "11", "01", "00", "01", "00", "01", "00", "11", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "11"),
463 => ("00", "00", "01", "00", "11", "00", "00", "00", "01", "11", "01", "01", "11", "11", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "11", "01", "01"),
464 => ("00", "00", "00", "00", "01", "11", "11", "00", "01", "01", "01", "11", "00", "00", "01", "11", "00", "00", "01", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00"),
465 => ("00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "11", "11", "11", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "11", "01"),
466 => ("00", "01", "01", "11", "00", "11", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "11", "11", "01", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "01"),
467 => ("01", "01", "01", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "11", "00", "11", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "00", "11", "11", "00", "00", "00"),
468 => ("01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01", "01", "11", "11", "01", "01", "11", "01", "00", "01", "00", "01", "11", "11", "00", "00", "00", "00", "00", "01"),
469 => ("00", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "00", "01", "11", "01", "00", "11", "01", "00", "01", "00", "11", "11", "00", "01", "01", "01", "11"),
470 => ("01", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "11", "00", "01", "00", "11", "11", "01", "11", "00", "11", "01", "01", "01", "01", "01", "01", "01"),
471 => ("00", "11", "01", "00", "01", "11", "01", "00", "00", "11", "00", "01", "01", "11", "11", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "01", "11", "00", "01", "01"),
472 => ("01", "11", "00", "11", "01", "00", "01", "00", "00", "00", "00", "11", "00", "11", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "11", "01", "11", "01", "01", "00", "00", "01"),
473 => ("01", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11", "11", "00", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11"),
474 => ("01", "11", "11", "01", "01", "01", "00", "01", "01", "01", "11", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00"),
475 => ("00", "00", "11", "01", "00", "00", "01", "11", "00", "00", "11", "11", "11", "00", "11", "01", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00"),
476 => ("01", "00", "00", "01", "00", "11", "11", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "11", "11", "00", "00", "00", "01", "01", "00"),
477 => ("00", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "11", "01", "00"),
478 => ("01", "01", "01", "11", "11", "00", "11", "00", "01", "01", "11", "01", "00", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "01", "11", "01", "01", "00", "01", "00"),
479 => ("00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "11", "00", "00", "11", "01", "01", "00", "01", "00", "11", "01", "00", "00", "01", "11", "11", "01"),
480 => ("00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "00", "01", "00", "00", "11", "01", "00", "11", "00", "11", "01", "11"),
481 => ("01", "01", "01", "00", "00", "00", "11", "11", "00", "11", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "11", "01", "01", "11"),
482 => ("01", "00", "00", "01", "01", "01", "11", "01", "00", "11", "00", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "11", "11", "01", "00", "00", "11"),
483 => ("00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "11", "11", "01", "11", "00", "01", "11", "00", "00", "11"),
484 => ("00", "11", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "01", "11", "01", "11", "00", "01", "01", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "11", "01", "01"),
485 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "11", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "11", "11", "01", "00", "00", "11", "01", "01", "00", "00"),
486 => ("01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "11", "01", "01", "01", "11", "01", "01", "01", "01", "00", "01", "00", "11", "11", "00", "00", "01", "01", "00"),
487 => ("00", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "11", "00", "11", "01", "01", "11", "11", "01", "00", "01", "01", "11", "01", "11"),
488 => ("00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "11", "01", "01", "11", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00"),
489 => ("01", "00", "01", "00", "01", "01", "11", "11", "11", "00", "00", "00", "11", "01", "00", "11", "01", "00", "01", "11", "01", "11", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00"),
490 => ("01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "11", "00", "01", "00", "01", "11", "11", "00", "11", "00"),
491 => ("00", "00", "01", "00", "00", "00", "11", "11", "00", "11", "00", "00", "00", "11", "00", "11", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00"),
492 => ("01", "01", "01", "11", "01", "11", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "11", "00", "11", "01", "01", "01", "00", "01", "01", "01"),
493 => ("01", "00", "11", "01", "01", "00", "00", "01", "01", "00", "11", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "01", "00", "11", "00", "11", "11", "00", "01", "00", "00", "11"),
494 => ("00", "11", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "11", "00", "01", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "00", "11", "00"),
495 => ("00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "11", "00", "00", "01", "00", "00", "11", "11", "01", "00", "01", "11", "00", "01", "01", "00", "01", "00", "01", "11"),
496 => ("00", "00", "01", "00", "01", "11", "01", "01", "11", "00", "00", "11", "11", "11", "00", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "01", "11", "00"),
497 => ("01", "11", "01", "01", "00", "11", "11", "01", "11", "01", "01", "01", "01", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00"),
498 => ("00", "11", "01", "11", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "11", "01", "11", "01"),
499 => ("00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "11", "11", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "11", "00", "11", "01", "01")),
(
0 => ("01", "00", "11", "00", "11", "11", "00", "01", "00", "11", "01", "11", "00", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01"),
1 => ("01", "01", "11", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "01", "01", "01", "00", "11", "00", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00"),
2 => ("00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "01", "00", "11", "00", "01", "11", "11", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "11"),
3 => ("00", "00", "11", "01", "01", "00", "01", "00", "11", "11", "11", "00", "01", "01", "00", "01", "01", "11", "11", "00", "00", "01", "11", "11", "01", "01", "00", "01", "01", "01", "00", "00"),
4 => ("00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "11", "00", "00", "11", "01", "11", "01", "00", "00", "11", "00", "11", "01", "00"),
5 => ("01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "01", "01", "01", "11", "00", "01", "11", "00", "00", "11", "01", "00", "01", "11", "01", "01", "01"),
6 => ("00", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "01", "11", "01", "11", "01", "01", "11", "01", "00"),
7 => ("01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "11", "11", "00", "00", "00", "01", "00", "11", "01", "01", "00", "11", "00", "00", "00", "11", "11", "00", "00"),
8 => ("01", "11", "11", "11", "00", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "11", "11", "00", "11", "00", "00", "00", "01", "00"),
9 => ("00", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "11", "11", "00", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "11", "11", "00"),
10 => ("01", "11", "01", "01", "01", "11", "01", "01", "00", "11", "00", "11", "00", "00", "11", "01", "00", "01", "01", "11", "11", "00", "01", "00", "01", "00", "01", "00", "01", "11", "01", "00"),
11 => ("01", "01", "00", "01", "11", "01", "01", "11", "01", "01", "11", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "11", "00", "11", "00", "00", "00"),
12 => ("01", "00", "00", "11", "11", "11", "01", "00", "11", "01", "11", "00", "01", "00", "11", "00", "00", "01", "11", "01", "00", "01", "00", "11", "00", "00", "00", "01", "00", "01", "00", "00"),
13 => ("01", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "11", "01", "11", "11", "01", "01", "11", "11", "01", "11", "00", "11", "01", "01", "01", "01", "00", "11", "01", "00", "01"),
14 => ("01", "01", "01", "01", "11", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "01", "11", "11", "01", "00", "01", "01", "11", "11", "00", "11", "00", "00", "01", "00", "01"),
15 => ("00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "11", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "11", "01", "11", "01"),
16 => ("01", "01", "01", "11", "01", "01", "01", "11", "01", "11", "01", "01", "01", "00", "01", "00", "11", "11", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "00", "00"),
17 => ("01", "00", "00", "00", "01", "00", "11", "11", "11", "11", "00", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00"),
18 => ("00", "11", "11", "00", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "11", "11", "00"),
19 => ("01", "11", "01", "00", "01", "01", "00", "00", "00", "11", "00", "00", "11", "11", "00", "00", "11", "11", "00", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00"),
20 => ("01", "11", "11", "01", "11", "01", "01", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "11", "01", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "11", "00", "01"),
21 => ("00", "11", "01", "01", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "11", "11", "01", "01", "00", "11", "01", "00", "01", "11", "01"),
22 => ("00", "01", "00", "11", "01", "00", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "11", "00", "01", "00", "11", "01", "00", "00", "11", "01", "01"),
23 => ("01", "01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "11", "00", "00", "11", "01", "01", "11", "00", "11", "01", "11", "01", "00", "00", "01", "00", "11", "00", "00", "01"),
24 => ("00", "00", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "00"),
25 => ("01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "11", "11", "11", "01", "11", "00", "00", "01", "11", "11", "00", "00", "00"),
26 => ("00", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "11", "11", "11", "01", "01", "01", "01", "00", "00", "11", "00", "11", "11", "00", "00", "01", "01", "00"),
27 => ("01", "00", "00", "00", "00", "01", "00", "11", "01", "01", "11", "01", "01", "00", "11", "00", "00", "00", "11", "11", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00"),
28 => ("00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "01", "01", "00", "01", "01", "11", "11", "11", "00", "11", "00", "11", "00", "11", "01", "00", "01", "00", "01", "01", "01", "01"),
29 => ("01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "11", "01", "00", "11", "11", "01"),
30 => ("01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "00", "00", "11", "01", "00", "11", "01", "00", "00", "01", "01", "11", "01", "00"),
31 => ("01", "01", "11", "11", "01", "00", "11", "00", "00", "01", "11", "00", "11", "01", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01"),
32 => ("00", "01", "11", "01", "11", "00", "00", "01", "11", "11", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "01", "11", "01", "11", "01", "00", "11", "00", "00", "01", "01"),
33 => ("00", "00", "00", "11", "00", "00", "01", "01", "11", "01", "11", "01", "01", "00", "01", "11", "01", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "00", "01"),
34 => ("01", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "00", "00", "00", "11", "01", "11", "11", "01", "01", "01", "01", "00", "11", "11", "01"),
35 => ("00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "11", "01", "11", "01", "01", "00", "11", "01", "11", "01", "00", "01", "00", "11", "00", "00", "11"),
36 => ("00", "00", "01", "00", "01", "01", "11", "00", "00", "11", "01", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "11", "01", "01", "01", "01", "00", "11", "01", "01", "00"),
37 => ("01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "01", "11", "11", "00", "11", "11"),
38 => ("01", "11", "01", "11", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "11", "00", "11", "11", "01", "01", "11", "00", "00", "00"),
39 => ("00", "00", "01", "00", "01", "00", "00", "01", "11", "11", "01", "11", "01", "01", "11", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00", "11", "00", "11", "01", "01", "00", "01"),
40 => ("00", "00", "11", "01", "11", "00", "01", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "01", "00", "00", "11", "00", "01", "11", "11", "00", "01", "01"),
41 => ("00", "01", "11", "01", "11", "01", "01", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "11", "01", "11", "01", "00", "01", "01", "11", "01"),
42 => ("01", "01", "11", "00", "01", "11", "01", "11", "00", "00", "00", "01", "00", "11", "11", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "01"),
43 => ("00", "00", "01", "01", "11", "00", "00", "00", "11", "11", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11", "11", "00", "00", "00", "11", "01", "00", "00", "11", "11"),
44 => ("01", "01", "00", "00", "11", "01", "01", "11", "00", "11", "01", "00", "00", "00", "01", "00", "11", "01", "11", "00", "00", "01", "00", "11", "11", "11", "00", "00", "01", "00", "00", "00"),
45 => ("00", "00", "11", "01", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11"),
46 => ("01", "01", "01", "00", "11", "00", "11", "11", "00", "11", "11", "11", "01", "00", "00", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "01", "11", "01", "01", "01", "00", "00"),
47 => ("01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "00", "11", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "11"),
48 => ("01", "00", "00", "01", "11", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "11", "11", "01"),
49 => ("00", "00", "01", "00", "11", "00", "01", "01", "00", "00", "11", "11", "01", "01", "00", "11", "01", "00", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "11", "11", "00"),
50 => ("01", "00", "00", "11", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "11", "11", "00", "11", "11", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "00", "00", "11"),
51 => ("00", "11", "00", "00", "11", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00"),
52 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "11", "11", "01", "01", "11", "01", "01", "00", "11", "11", "01", "01", "01", "01", "00", "11"),
53 => ("00", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "01", "01", "01", "00", "11", "01", "01", "01", "00"),
54 => ("00", "00", "00", "01", "00", "11", "11", "01", "00", "01", "00", "00", "11", "11", "01", "00", "00", "00", "11", "00", "11", "00", "01", "00", "01", "11", "01", "01", "01", "00", "11", "01"),
55 => ("00", "00", "01", "00", "11", "01", "11", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "00", "11", "01", "11", "00", "11", "01", "01", "00", "01", "00", "01"),
56 => ("01", "01", "00", "01", "11", "01", "00", "00", "11", "01", "00", "11", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "00"),
57 => ("00", "01", "11", "00", "00", "01", "01", "01", "11", "11", "11", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "00", "00"),
58 => ("01", "00", "11", "11", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "01", "11", "01", "01", "01", "01", "00"),
59 => ("00", "01", "01", "01", "00", "01", "11", "00", "01", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "11", "11", "11", "01", "01", "11", "00", "00", "00"),
60 => ("00", "00", "01", "01", "01", "11", "00", "11", "01", "11", "11", "01", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01"),
61 => ("00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "11", "00", "01", "01", "11", "01", "00", "11", "01", "01", "00", "01", "00", "11", "00", "01", "01"),
62 => ("01", "11", "01", "00", "00", "00", "11", "00", "11", "01", "00", "00", "11", "01", "11", "01", "11", "00", "01", "01", "11", "00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "00"),
63 => ("01", "01", "11", "01", "00", "01", "00", "00", "01", "11", "11", "01", "11", "01", "11", "01", "01", "00", "00", "01", "00", "11", "11", "00", "11", "01", "01", "01", "01", "01", "00", "00"),
64 => ("00", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "11", "01", "11", "01", "00", "11", "00", "01", "01", "11", "01", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01"),
65 => ("00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "11", "01", "00", "11", "00", "00", "01", "00", "01", "00", "11", "01", "11", "00", "00", "11", "01", "11", "01", "00", "01"),
66 => ("00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "11", "00", "01", "01", "00", "01"),
67 => ("00", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "11", "11", "11", "01", "11", "00", "11", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01"),
68 => ("00", "01", "01", "01", "11", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "11", "11", "00", "01", "11", "11", "11", "01", "11", "00", "00", "01", "01", "01", "00"),
69 => ("00", "11", "01", "00", "00", "01", "00", "01", "00", "00", "11", "11", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "00", "00", "11", "00", "11", "00", "01", "01", "01", "01"),
70 => ("00", "11", "01", "11", "11", "01", "01", "11", "01", "00", "01", "01", "11", "01", "11", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00"),
71 => ("01", "00", "01", "01", "01", "11", "01", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "11", "11", "11", "00", "01", "00", "00", "01", "01"),
72 => ("00", "11", "00", "00", "01", "00", "01", "00", "01", "01", "01", "00", "11", "01", "01", "00", "00", "01", "00", "11", "01", "11", "11", "01", "01", "01", "01", "01", "11", "11", "00", "01"),
73 => ("00", "01", "11", "00", "11", "11", "00", "00", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "00", "11", "01", "00", "00", "11", "00", "01", "01", "00", "11", "01", "01", "01"),
74 => ("00", "00", "01", "01", "00", "11", "11", "11", "01", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "00", "11", "11", "01", "11", "00", "01", "00", "00"),
75 => ("01", "11", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "00", "11", "00", "01", "00", "00", "00", "01", "00"),
76 => ("01", "01", "11", "01", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "01", "11", "11", "00"),
77 => ("00", "11", "00", "01", "01", "00", "11", "11", "11", "00", "01", "01", "00", "01", "01", "01", "11", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "00", "11", "00", "01", "00"),
78 => ("01", "00", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "11", "00", "00", "11", "11", "11", "00", "01", "11", "11", "00", "01", "11", "01", "00", "00", "00", "00", "00"),
79 => ("00", "00", "11", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "00", "11"),
80 => ("01", "00", "00", "11", "01", "01", "11", "00", "00", "00", "00", "01", "00", "11", "01", "11", "00", "01", "11", "01", "00", "00", "01", "00", "00", "11", "00", "01", "11", "00", "00", "01"),
81 => ("01", "00", "00", "11", "01", "11", "01", "00", "00", "11", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "11", "00", "01", "00", "01", "11", "01", "01"),
82 => ("00", "01", "01", "00", "11", "00", "01", "11", "00", "01", "01", "00", "11", "00", "11", "00", "00", "00", "01", "01", "11", "01", "11", "00", "01", "01", "00", "00", "11", "00", "00", "01"),
83 => ("00", "00", "11", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "11", "00", "00", "01", "00", "01", "11", "00", "00", "00", "11", "01", "11"),
84 => ("00", "11", "11", "01", "11", "00", "01", "00", "00", "01", "11", "11", "01", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "01", "01", "00", "11", "00", "11", "11", "00", "01"),
85 => ("00", "01", "01", "01", "11", "00", "00", "01", "01", "11", "11", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "11", "01", "01", "01", "11"),
86 => ("01", "01", "01", "11", "00", "01", "01", "01", "11", "01", "11", "11", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00"),
87 => ("01", "01", "01", "01", "00", "11", "00", "00", "11", "00", "11", "00", "00", "00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "11"),
88 => ("01", "01", "00", "11", "00", "01", "01", "00", "11", "11", "00", "11", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01"),
89 => ("00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "00", "00", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "11", "01"),
90 => ("00", "11", "00", "01", "11", "11", "01", "11", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "11", "00", "11", "01", "01", "00", "01", "01", "00"),
91 => ("00", "01", "00", "00", "00", "00", "11", "11", "11", "01", "00", "00", "11", "00", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "11", "00", "00", "01"),
92 => ("01", "01", "00", "01", "11", "11", "01", "11", "01", "01", "01", "00", "00", "11", "00", "01", "01", "11", "00", "00", "01", "01", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01"),
93 => ("00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "00", "11", "11", "11", "11", "11", "01", "01", "11", "01", "01", "01", "01", "11", "00", "00"),
94 => ("00", "01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "00", "00", "01", "11", "11", "11", "01", "01", "00", "01", "00", "00", "00", "11", "11", "01", "01", "11", "01", "00"),
95 => ("00", "01", "00", "00", "01", "00", "01", "11", "11", "11", "01", "00", "11", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "11", "01", "11", "01", "01", "01", "11", "01", "01"),
96 => ("00", "00", "00", "11", "11", "11", "01", "01", "01", "00", "11", "11", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "00"),
97 => ("00", "01", "00", "01", "11", "11", "01", "00", "01", "00", "11", "00", "00", "11", "00", "01", "00", "00", "01", "00", "01", "11", "01", "01", "01", "11", "01", "01", "00", "11", "01", "01"),
98 => ("00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "11", "11", "00", "01", "00", "00", "00", "00", "01", "11", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "11"),
99 => ("00", "11", "01", "00", "00", "01", "00", "11", "00", "01", "01", "11", "01", "01", "01", "01", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "11", "00", "11", "01"),
100 => ("00", "00", "11", "11", "01", "00", "01", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "11", "11", "00", "01", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "00"),
101 => ("00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "11", "11", "11", "00", "11"),
102 => ("01", "00", "11", "00", "11", "00", "00", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "11", "00", "11", "11"),
103 => ("01", "00", "00", "11", "00", "01", "11", "00", "01", "00", "00", "01", "11", "00", "00", "01", "00", "01", "01", "00", "11", "11", "11", "11", "01", "01", "00", "11", "01", "01", "01", "01"),
104 => ("01", "01", "00", "00", "01", "01", "11", "11", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "11", "11", "00", "01", "01", "00", "00", "00", "01", "11", "11", "00", "00", "01"),
105 => ("00", "01", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "00", "01", "00", "01", "11", "00", "00", "00", "11", "00", "01", "01", "11", "01"),
106 => ("00", "00", "01", "01", "00", "11", "00", "00", "11", "00", "01", "11", "11", "01", "01", "00", "01", "11", "00", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01"),
107 => ("01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "11", "11", "01", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "11", "01", "00", "01", "01", "01", "11", "00", "00"),
108 => ("01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "11", "01", "11", "00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "11", "01", "00", "01"),
109 => ("00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "01", "00", "01", "11", "01", "01", "01", "01", "00", "11", "00", "00", "00", "11", "11", "00", "00", "00", "11"),
110 => ("01", "00", "00", "00", "00", "00", "11", "00", "01", "00", "11", "11", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "01", "01", "00"),
111 => ("01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "01", "00", "00", "11", "01", "00", "01", "01", "11", "11", "00", "01", "00", "00", "11", "11", "01", "01"),
112 => ("01", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "11", "11", "01", "11", "00", "01", "11", "00", "01", "01", "11", "00"),
113 => ("01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "01", "11"),
114 => ("00", "01", "00", "00", "11", "01", "00", "00", "01", "00", "01", "11", "01", "11", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "00", "11", "11", "01", "00", "01", "00", "00"),
115 => ("01", "11", "01", "00", "11", "01", "00", "01", "11", "00", "11", "11", "00", "00", "01", "01", "00", "01", "00", "01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "01", "00", "11"),
116 => ("01", "01", "00", "11", "01", "00", "11", "00", "01", "11", "00", "11", "11", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "00", "00", "00", "00"),
117 => ("01", "00", "11", "00", "01", "11", "01", "01", "01", "01", "01", "11", "00", "11", "00", "11", "01", "01", "00", "00", "01", "11", "00", "01", "11", "00", "00", "01", "11", "01", "00", "00"),
118 => ("00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "11", "01", "01", "01", "00", "00", "01", "11", "11"),
119 => ("01", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "00", "01", "11", "00", "11", "01", "00", "01", "00", "00", "11", "11", "01", "11", "00", "01", "01"),
120 => ("00", "01", "11", "11", "01", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "00"),
121 => ("01", "01", "01", "11", "01", "01", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "11", "01", "01", "11", "11", "11", "00", "01", "01", "01", "11", "01"),
122 => ("01", "11", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "11", "11", "11", "00", "00", "00", "11"),
123 => ("01", "00", "01", "00", "11", "01", "00", "11", "11", "00", "01", "00", "00", "11", "01", "00", "11", "00", "11", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11"),
124 => ("00", "11", "11", "01", "11", "11", "01", "00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01"),
125 => ("01", "11", "01", "11", "11", "11", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "11", "00", "00", "01", "11", "01", "00", "00", "11", "00", "00", "01", "00", "01", "00", "01"),
126 => ("00", "01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "11", "11", "00", "00", "11", "00", "11", "01", "11", "01", "01", "00", "11", "11"),
127 => ("00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "00", "11", "00", "01", "11", "00", "11", "01", "01", "11", "00", "00", "00", "01"),
128 => ("01", "00", "00", "11", "01", "11", "01", "11", "01", "01", "01", "01", "11", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "00", "00", "01", "00", "11", "11", "00"),
129 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "00", "00", "11", "01", "01", "00", "11", "00", "11", "01", "00", "01", "11", "11", "00", "11", "01", "11"),
130 => ("01", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "01", "11", "01", "01", "11", "00", "01", "11", "01", "01", "01", "11", "01", "00", "11"),
131 => ("01", "11", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "11", "01", "01", "01", "11", "01", "01", "00", "11"),
132 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "01", "01", "01", "11", "01", "01", "11", "11", "00", "11", "00"),
133 => ("01", "00", "01", "00", "11", "11", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "11", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01"),
134 => ("01", "01", "00", "00", "11", "00", "00", "01", "00", "11", "11", "01", "01", "00", "11", "01", "00", "00", "11", "00", "01", "01", "00", "01", "00", "00", "00", "11", "11", "11", "00", "00"),
135 => ("01", "11", "01", "00", "11", "11", "01", "11", "00", "00", "00", "00", "00", "00", "01", "00", "11", "11", "01", "11", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00"),
136 => ("00", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "11", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "11", "00", "00", "00", "11", "11", "11", "00", "00"),
137 => ("01", "00", "01", "11", "00", "00", "11", "00", "01", "11", "00", "11", "01", "11", "01", "01", "11", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "11", "00", "01", "00", "01"),
138 => ("00", "00", "00", "11", "01", "00", "00", "01", "11", "11", "01", "01", "01", "11", "11", "01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "11"),
139 => ("01", "00", "11", "11", "01", "01", "00", "01", "01", "00", "11", "00", "11", "11", "01", "11", "00", "00", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "11", "01"),
140 => ("01", "01", "00", "00", "11", "00", "00", "00", "11", "00", "11", "00", "11", "11", "01", "01", "11", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "00"),
141 => ("01", "00", "00", "11", "00", "11", "11", "00", "11", "00", "01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "11", "00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "00"),
142 => ("01", "11", "01", "01", "00", "11", "00", "11", "00", "01", "00", "11", "00", "11", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00", "11", "01", "00", "00", "00", "01", "00", "00"),
143 => ("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "11", "11", "11", "11", "11", "11", "00", "01", "00", "00"),
144 => ("01", "11", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "11", "11", "00", "01", "00", "11", "00", "01", "11", "00", "11", "00", "00", "01", "00", "00", "00", "11", "01"),
145 => ("01", "00", "11", "00", "01", "11", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "11", "01", "00", "11", "00", "01", "01", "01", "01", "01", "01", "11", "01", "11", "00", "01"),
146 => ("01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "01", "01", "01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "11", "00"),
147 => ("01", "01", "11", "11", "00", "00", "01", "01", "00", "11", "00", "00", "11", "01", "00", "00", "00", "01", "01", "11", "01", "00", "11", "01", "00", "00", "11", "00", "00", "11", "01", "01"),
148 => ("01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "01", "01", "11", "00", "11", "11", "01", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "11", "11", "00", "00", "11"),
149 => ("01", "01", "01", "00", "01", "01", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "11", "11", "11", "00", "00", "00", "01", "11", "01", "00", "11", "00", "11", "00", "11", "01"),
150 => ("00", "00", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "11", "00", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "11"),
151 => ("00", "01", "01", "01", "11", "01", "00", "11", "01", "01", "00", "00", "00", "11", "11", "01", "11", "00", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "00", "00", "11", "01"),
152 => ("00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "00", "01", "01", "11", "00", "01", "11", "00", "01", "00", "11", "01", "11", "01", "01", "11", "11", "01", "00", "01", "00"),
153 => ("01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "11", "11", "01", "00", "01", "00", "00", "00", "00", "11", "00", "11", "00", "00", "01", "11", "01", "11"),
154 => ("00", "00", "11", "01", "01", "01", "01", "11", "11", "11", "01", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00"),
155 => ("01", "11", "11", "00", "01", "00", "11", "01", "11", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "00"),
156 => ("01", "01", "00", "00", "11", "11", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01"),
157 => ("00", "00", "11", "11", "01", "11", "00", "00", "00", "01", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "11", "00", "00", "11", "01", "00", "11", "11"),
158 => ("01", "11", "00", "01", "11", "01", "11", "00", "01", "01", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "01", "01", "00"),
159 => ("00", "11", "00", "01", "11", "11", "00", "00", "00", "01", "11", "11", "00", "00", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00"),
160 => ("00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "11", "00", "11", "01", "00", "01", "01", "00", "01", "11", "01", "01", "00", "01", "00", "11", "00", "00", "00", "11", "01", "11"),
161 => ("01", "11", "01", "01", "00", "11", "11", "00", "00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "01"),
162 => ("01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "11", "11", "01", "00", "11", "11", "00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "01", "00"),
163 => ("01", "11", "00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "11", "01", "00", "01", "00", "11", "00", "01", "11", "01", "11", "01", "00", "00", "00", "01", "11", "01", "01"),
164 => ("00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "11", "01", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "00", "01", "11", "00", "00", "11", "01", "11", "01", "00"),
165 => ("01", "01", "01", "00", "01", "11", "11", "01", "01", "11", "00", "11", "01", "00", "00", "01", "01", "01", "11", "11", "00", "00", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00"),
166 => ("01", "01", "01", "11", "11", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "11", "01", "00", "00", "11"),
167 => ("01", "00", "00", "00", "11", "00", "11", "00", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "00", "11", "11", "11", "00", "01", "00"),
168 => ("00", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "11", "01", "01", "00", "01", "11", "11", "01", "11", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01"),
169 => ("01", "01", "11", "01", "01", "01", "00", "11", "01", "00", "01", "11", "01", "11", "00", "00", "01", "00", "11", "01", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01"),
170 => ("01", "01", "00", "00", "11", "00", "00", "01", "11", "11", "11", "00", "00", "01", "01", "00", "00", "01", "11", "01", "01", "11", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00"),
171 => ("01", "00", "11", "11", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "01", "11", "00", "01", "01", "01", "00", "00", "00", "11", "00", "11", "00", "01", "00", "11", "00", "01"),
172 => ("01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "11", "01", "00", "00", "11", "01", "11", "00", "00", "00", "11", "00", "01", "01", "11", "11", "00", "01", "01", "11", "01", "01"),
173 => ("01", "00", "01", "01", "11", "11", "01", "01", "01", "01", "01", "01", "00", "11", "11", "11", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "11"),
174 => ("01", "11", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "11", "11", "01", "00", "00", "00", "00", "11", "00", "01", "00", "11", "11", "11", "00", "11", "01", "00"),
175 => ("01", "11", "00", "01", "11", "11", "01", "01", "00", "00", "01", "00", "01", "00", "11", "01", "11", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "01"),
176 => ("00", "01", "00", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "11", "11", "11", "00", "11"),
177 => ("00", "01", "01", "01", "00", "00", "11", "11", "01", "11", "00", "01", "00", "11", "01", "01", "01", "01", "01", "11", "11", "01", "11", "11", "01", "00", "01", "01", "01", "00", "00", "00"),
178 => ("00", "11", "01", "00", "11", "01", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "11", "11", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "00", "11", "00"),
179 => ("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "11", "01", "11", "11", "01", "00", "11", "00", "00", "00", "11", "01", "00", "01", "00", "00", "00", "11", "01", "11"),
180 => ("01", "11", "01", "01", "01", "01", "00", "01", "00", "11", "11", "01", "11", "00", "01", "01", "11", "11", "00", "01", "01", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01"),
181 => ("01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "11", "01", "11", "00", "00", "01"),
182 => ("00", "11", "00", "00", "01", "11", "00", "01", "01", "00", "01", "00", "11", "01", "00", "11", "00", "01", "01", "11", "00", "00", "01", "01", "11", "01", "00", "11", "01", "01", "11", "00"),
183 => ("00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "11", "11", "11", "00", "01", "00", "01", "11"),
184 => ("01", "11", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "00", "01", "00", "00", "01", "00", "11", "01", "01", "01", "11", "00", "01", "01", "00", "11", "00"),
185 => ("00", "00", "00", "01", "11", "00", "01", "00", "11", "11", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "01", "11", "00", "01", "00"),
186 => ("01", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01", "11", "00", "00", "11", "00", "11", "11", "00", "11", "00", "01", "01", "11", "00", "01", "01", "01", "01"),
187 => ("00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "01", "11", "00", "00", "11", "00"),
188 => ("00", "00", "01", "00", "01", "11", "01", "01", "00", "01", "11", "01", "00", "11", "11", "01", "00", "00", "11", "01", "00", "11", "00", "11", "01", "00", "01", "11", "01", "00", "01", "00"),
189 => ("01", "00", "00", "00", "01", "11", "11", "00", "11", "11", "00", "11", "01", "11", "00", "01", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00"),
190 => ("01", "11", "11", "11", "01", "01", "11", "01", "01", "11", "00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "11"),
191 => ("01", "11", "01", "01", "11", "01", "01", "00", "01", "00", "11", "01", "11", "11", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "00", "01", "01", "11", "00", "00"),
192 => ("01", "01", "11", "01", "11", "00", "00", "00", "01", "11", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "01", "11", "11", "01"),
193 => ("01", "01", "00", "01", "11", "00", "11", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "00", "11", "11", "01", "00", "01", "00", "01", "00", "00", "00", "00", "01", "01", "11"),
194 => ("00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "01", "11", "00", "01", "01", "11", "00", "01", "11", "11", "00", "01", "00", "01", "01", "11", "00", "11", "01", "00", "00"),
195 => ("01", "01", "11", "00", "00", "01", "01", "11", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "01", "11", "01", "00", "11", "00", "11", "00", "01", "11", "00", "00"),
196 => ("01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "01", "01", "01", "11", "00", "11", "11", "11", "00", "11", "00", "01", "00", "00", "01"),
197 => ("01", "01", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "00", "00", "01", "00", "00", "11", "00", "11", "01", "01", "01", "00", "00", "01", "01", "11", "11", "01", "01"),
198 => ("00", "00", "01", "01", "01", "11", "11", "00", "00", "01", "11", "01", "00", "11", "00", "00", "01", "00", "01", "01", "11", "11", "01", "11", "01", "01", "00", "00", "11", "01", "01", "01"),
199 => ("00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "11", "01", "00", "00", "01", "01", "11", "00", "11", "00", "11", "11", "00", "01", "00"),
200 => ("00", "00", "01", "01", "00", "11", "00", "01", "01", "00", "11", "00", "00", "11", "00", "00", "01", "01", "01", "11", "11", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "11"),
201 => ("00", "01", "00", "01", "11", "01", "00", "11", "00", "00", "01", "01", "01", "00", "00", "00", "11", "11", "00", "01", "00", "01", "11", "01", "01", "01", "11", "01", "01", "11", "01", "01"),
202 => ("01", "01", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "01", "11", "11", "00", "01", "11", "11", "11", "00", "00"),
203 => ("01", "01", "11", "01", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "00", "01", "00", "01", "11", "01", "00", "01", "11", "01", "01", "11", "01", "01"),
204 => ("00", "00", "01", "00", "01", "11", "01", "11", "11", "00", "00", "00", "00", "11", "11", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01"),
205 => ("00", "01", "00", "11", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "01", "00", "11", "01", "11", "11", "01", "00", "01", "11", "00", "01"),
206 => ("00", "01", "00", "01", "00", "00", "01", "01", "00", "01", "00", "01", "00", "01", "11", "11", "00", "11", "00", "01", "01", "11", "00", "11", "01", "11", "00", "11", "00", "00", "01", "01"),
207 => ("00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "11", "00", "01", "11", "11", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "11", "01", "11", "01", "01", "11"),
208 => ("01", "11", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "01", "11", "01", "11", "00", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11"),
209 => ("00", "01", "11", "11", "01", "00", "11", "01", "11", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00"),
210 => ("00", "01", "00", "11", "00", "01", "00", "00", "11", "00", "01", "11", "01", "00", "01", "01", "11", "11", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00"),
211 => ("01", "01", "00", "00", "11", "01", "11", "01", "01", "00", "00", "01", "00", "11", "00", "00", "00", "11", "00", "00", "00", "11", "01", "01", "11", "11", "00", "00", "00", "01", "00", "01"),
212 => ("00", "01", "01", "00", "00", "11", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "01", "00", "01", "01", "11", "11", "11", "11", "01", "00", "01", "11"),
213 => ("00", "00", "11", "01", "01", "11", "00", "00", "00", "00", "00", "11", "01", "01", "00", "00", "01", "11", "00", "00", "01", "11", "01", "11", "11", "00", "00", "00", "01", "00", "00", "11"),
214 => ("01", "00", "01", "00", "01", "00", "11", "11", "11", "01", "00", "01", "00", "11", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "00", "01", "00"),
215 => ("00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "11", "01", "01", "00", "01", "01", "01", "00", "11", "00", "11", "00", "11", "01", "11", "11", "01", "00", "00"),
216 => ("00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "00", "01", "11", "11", "00", "01", "01", "11", "11", "11"),
217 => ("01", "11", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "01", "11", "11", "00", "11", "00", "00", "11", "00", "11"),
218 => ("00", "11", "01", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "11", "11", "00", "01", "00", "11", "01", "01", "00", "11", "00", "01", "01", "01", "00", "01", "01", "11"),
219 => ("01", "01", "01", "11", "00", "00", "00", "01", "00", "01", "01", "11", "00", "11", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "11", "01", "11", "11", "00", "01"),
220 => ("00", "00", "01", "00", "01", "00", "01", "01", "00", "11", "11", "01", "11", "11", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "11", "01", "11", "11", "01", "00", "00", "01"),
221 => ("01", "01", "01", "00", "00", "00", "00", "00", "11", "01", "11", "11", "11", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "11", "01", "00", "00", "01", "01", "00", "00", "11"),
222 => ("01", "11", "00", "01", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "00", "11", "00", "11", "00", "01", "01", "11", "11", "00", "00"),
223 => ("00", "11", "00", "00", "01", "00", "01", "11", "01", "11", "01", "01", "01", "11", "01", "01", "00", "11", "00", "01", "00", "01", "00", "00", "00", "11", "00", "00", "00", "01", "11", "11"),
224 => ("01", "00", "01", "00", "00", "11", "01", "01", "01", "11", "01", "00", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "11", "01", "00", "00", "01", "11", "01", "11", "01"),
225 => ("01", "11", "11", "01", "11", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "00", "01", "01", "01", "01", "00", "00", "11", "11", "00", "01", "01", "11", "11", "00"),
226 => ("00", "11", "00", "00", "11", "00", "11", "00", "01", "00", "00", "11", "01", "11", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "01", "11", "01"),
227 => ("00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "11", "00", "00"),
228 => ("00", "00", "11", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "11", "00", "01", "00", "11", "01", "01"),
229 => ("00", "01", "11", "01", "00", "11", "11", "00", "00", "01", "01", "11", "01", "00", "00", "11", "11", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11"),
230 => ("01", "01", "00", "11", "01", "01", "11", "00", "01", "00", "00", "00", "11", "01", "01", "01", "00", "00", "01", "00", "01", "11", "11", "11", "01", "00", "00", "01", "00", "00", "11", "11"),
231 => ("00", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "11", "11", "01", "11", "00", "11", "01", "11", "01", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "01", "11"),
232 => ("00", "00", "00", "00", "00", "11", "00", "01", "01", "01", "11", "11", "11", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "11", "00", "00", "00", "11", "01", "00", "00"),
233 => ("01", "01", "00", "11", "01", "01", "11", "01", "00", "01", "01", "11", "01", "11", "01", "11", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "11", "00", "01"),
234 => ("00", "00", "11", "00", "00", "01", "01", "11", "00", "00", "01", "11", "01", "01", "01", "01", "11", "11", "00", "01", "00", "00", "00", "01", "11", "01", "00", "11", "00", "00", "00", "01"),
235 => ("01", "11", "01", "01", "00", "00", "00", "11", "11", "00", "01", "11", "01", "00", "01", "11", "11", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01", "01", "11", "00"),
236 => ("01", "00", "11", "00", "00", "00", "00", "11", "00", "11", "01", "11", "11", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00", "01", "11", "01", "01", "01"),
237 => ("01", "00", "11", "01", "11", "01", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "00", "11", "01", "01", "00", "01", "00", "00", "11", "01", "00"),
238 => ("00", "01", "01", "01", "11", "11", "11", "01", "01", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01"),
239 => ("00", "00", "00", "00", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "11", "00", "11", "01", "00", "00", "00", "00", "01", "11", "01", "01", "11", "11", "00", "00"),
240 => ("00", "00", "11", "00", "01", "11", "00", "11", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01"),
241 => ("01", "01", "00", "01", "11", "00", "00", "01", "11", "00", "00", "01", "01", "00", "00", "11", "00", "01", "11", "01", "00", "01", "01", "11", "00", "01", "11", "00", "01", "01", "00", "11"),
242 => ("00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "11", "01", "01", "11", "11", "01", "00", "00", "00", "11", "00", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00"),
243 => ("00", "01", "11", "11", "00", "11", "01", "01", "01", "11", "01", "00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "01", "00", "00"),
244 => ("01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "01", "11", "00", "00", "00", "11", "11", "00", "01", "11", "01", "01", "00", "00", "01", "11", "00", "00", "00"),
245 => ("01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "11", "01", "11", "01", "11", "00", "00", "11", "11", "00", "00", "01", "00", "11", "11", "00"),
246 => ("01", "01", "11", "01", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "11", "11", "01", "01", "00", "11", "00", "00"),
247 => ("00", "11", "01", "00", "00", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "11", "01", "11"),
248 => ("01", "11", "01", "00", "01", "00", "11", "01", "11", "01", "01", "11", "11", "11", "01", "01", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00"),
249 => ("00", "01", "00", "11", "01", "01", "11", "01", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "11", "00", "11", "01"),
250 => ("01", "11", "01", "00", "01", "01", "00", "01", "01", "01", "11", "11", "11", "01", "00", "00", "00", "00", "00", "01", "00", "11", "00", "11", "01", "01", "01", "11", "01", "01", "01", "01"),
251 => ("01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "11", "11", "11", "01", "01", "00", "11", "11", "00", "01", "00", "01", "00", "11"),
252 => ("00", "01", "01", "00", "00", "01", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "01", "11", "11", "01", "11", "01", "01", "11", "01", "00", "00", "01", "00", "11", "00", "00"),
253 => ("01", "11", "00", "00", "11", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "11", "11", "01", "11", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00"),
254 => ("00", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "00", "11", "01", "00", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "11", "00", "11", "00", "01", "01", "00"),
255 => ("01", "01", "00", "01", "00", "11", "11", "01", "01", "01", "00", "11", "00", "00", "00", "01", "11", "11", "00", "01", "01", "11", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01"),
256 => ("01", "00", "01", "01", "00", "01", "11", "00", "11", "00", "01", "00", "11", "01", "00", "11", "01", "00", "01", "01", "00", "11", "00", "00", "00", "00", "11", "01", "11", "01", "00", "01"),
257 => ("01", "00", "00", "01", "01", "00", "00", "01", "11", "11", "00", "11", "11", "00", "00", "11", "00", "00", "01", "11", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "00"),
258 => ("01", "01", "11", "11", "11", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "01", "00", "11", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "11", "01", "01", "11"),
259 => ("01", "00", "01", "01", "01", "11", "01", "11", "11", "00", "01", "01", "00", "11", "01", "00", "11", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "01", "00", "11", "11"),
260 => ("00", "11", "11", "01", "01", "11", "00", "01", "11", "01", "01", "01", "00", "11", "00", "00", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "00", "11", "01", "11"),
261 => ("00", "01", "11", "00", "01", "00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11", "11", "00", "00", "00"),
262 => ("00", "11", "01", "01", "01", "11", "01", "11", "01", "00", "11", "11", "01", "01", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "11", "01", "01", "01"),
263 => ("01", "11", "00", "01", "01", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "11", "00", "00", "01", "00", "01", "11", "00", "11", "11", "01", "01", "01", "00", "01", "11"),
264 => ("01", "11", "11", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "00", "01", "00", "00", "01", "01", "01", "01", "11", "00", "01", "11", "01", "00", "01", "11", "00", "01", "00"),
265 => ("01", "00", "00", "01", "00", "11", "01", "00", "11", "01", "01", "01", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "11", "11", "01", "01", "11", "01"),
266 => ("01", "01", "00", "01", "11", "11", "00", "01", "00", "01", "11", "01", "11", "01", "01", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "00", "01"),
267 => ("00", "01", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "11", "00", "01", "01", "01", "01", "01", "11", "00", "11", "11", "01", "11", "01", "01", "01", "01", "00", "00", "00"),
268 => ("00", "00", "00", "00", "00", "00", "01", "11", "01", "11", "11", "01", "01", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "11", "00", "00", "01", "11", "11", "01", "11", "00"),
269 => ("00", "00", "01", "11", "11", "11", "00", "00", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "11", "00", "01", "01"),
270 => ("00", "00", "01", "11", "01", "00", "01", "01", "11", "00", "01", "00", "00", "01", "01", "00", "01", "01", "00", "11", "11", "01", "00", "11", "00", "01", "01", "00", "00", "11", "00", "01"),
271 => ("01", "00", "11", "11", "00", "11", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "00", "01", "11", "01", "11", "01", "11", "11", "01"),
272 => ("00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "11", "00", "11", "00", "11", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "11", "01", "00"),
273 => ("00", "00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "11", "11", "01", "00", "00", "00", "11", "01", "01", "01", "01", "11", "01", "11", "11", "00", "01", "00"),
274 => ("01", "11", "01", "01", "11", "00", "01", "00", "11", "00", "01", "11", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "11", "01", "01", "11", "11", "01", "00"),
275 => ("01", "00", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "11", "11", "11", "00", "00", "11", "00", "11", "11"),
276 => ("00", "01", "11", "11", "01", "11", "11", "01", "01", "01", "00", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "11", "01", "11", "00", "01", "01"),
277 => ("01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "11", "01", "01", "00", "11", "01", "01", "00", "11", "00"),
278 => ("00", "01", "00", "11", "00", "00", "00", "01", "01", "11", "01", "11", "00", "00", "00", "11", "01", "01", "11", "01", "00", "01", "11", "01", "11", "00", "00", "01", "11", "01", "00", "00"),
279 => ("01", "11", "00", "01", "01", "11", "11", "01", "01", "11", "00", "11", "01", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "00", "01", "00"),
280 => ("00", "00", "01", "00", "11", "00", "01", "01", "00", "11", "01", "01", "01", "11", "01", "01", "01", "11", "01", "01", "11", "01", "01", "00", "01", "11", "01", "00", "01", "01", "01", "00"),
281 => ("01", "00", "00", "01", "01", "11", "11", "00", "00", "11", "00", "01", "00", "11", "11", "01", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "11", "01"),
282 => ("01", "01", "00", "00", "00", "11", "11", "01", "01", "01", "11", "00", "11", "01", "01", "00", "00", "00", "00", "00", "01", "01", "11", "01", "00", "11", "11", "01", "11", "01", "01", "00"),
283 => ("01", "01", "11", "11", "01", "01", "11", "00", "01", "01", "01", "11", "01", "00", "00", "11", "11", "11", "01", "00", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "00", "01"),
284 => ("01", "01", "11", "01", "00", "01", "01", "11", "11", "00", "11", "01", "01", "00", "11", "11", "00", "01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "00", "11", "00", "00"),
285 => ("00", "01", "00", "01", "00", "11", "01", "00", "00", "00", "11", "00", "00", "00", "11", "00", "00", "11", "00", "01", "01", "01", "11", "01", "00", "11", "11", "01", "00", "00", "00", "01"),
286 => ("01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00", "11", "00", "01", "00", "01", "01", "01", "11", "01", "11", "11", "01", "01", "01", "00", "00", "00", "11"),
287 => ("01", "11", "00", "00", "00", "11", "00", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "11", "01"),
288 => ("00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "00", "00", "00", "01", "01", "01", "00", "11", "11", "01", "11", "11", "11", "00", "00", "00", "01", "00"),
289 => ("00", "00", "11", "00", "00", "01", "11", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "00", "00", "00", "00", "11"),
290 => ("00", "01", "11", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "00", "01", "01", "11", "01", "11", "00", "01", "00", "01", "11", "01", "11", "00"),
291 => ("00", "00", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "11", "00", "01", "00", "11", "00", "11", "11", "01", "00", "11", "00", "01", "11"),
292 => ("00", "11", "01", "01", "01", "01", "01", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "11", "11", "00", "01", "01", "00", "00", "00", "00", "11", "00", "11", "01", "00", "00"),
293 => ("00", "11", "01", "01", "01", "11", "00", "00", "11", "01", "11", "11", "01", "00", "11", "01", "00", "00", "00", "00", "11", "01", "00", "00", "01", "11", "00", "01", "01", "00", "01", "01"),
294 => ("00", "00", "01", "11", "01", "00", "11", "00", "00", "00", "01", "00", "01", "11", "11", "11", "11", "00", "00", "01", "01", "00", "01", "01", "11", "01", "01", "11", "01", "01", "01", "01"),
295 => ("00", "00", "11", "01", "00", "01", "00", "01", "00", "11", "01", "11", "00", "00", "01", "11", "01", "11", "01", "00", "01", "01", "00", "11", "00", "01", "01", "01", "01", "00", "11", "01"),
296 => ("01", "01", "11", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00", "00", "00", "11", "00", "00", "00", "11", "01", "11"),
297 => ("01", "01", "01", "00", "01", "00", "01", "01", "11", "01", "00", "00", "11", "00", "11", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "11", "00", "01", "01", "11"),
298 => ("00", "00", "11", "11", "00", "00", "01", "00", "00", "01", "01", "01", "01", "00", "01", "00", "00", "01", "11", "01", "00", "11", "11", "01", "00", "11", "00", "11", "00", "11", "00", "01"),
299 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "01", "11", "00", "01", "11", "00", "00", "11", "00", "11", "01", "00", "11", "00", "00", "11", "01", "00", "01", "00", "11"),
300 => ("01", "00", "11", "11", "01", "00", "01", "11", "01", "00", "00", "00", "01", "11", "11", "01", "00", "01", "01", "11", "01", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00", "00"),
301 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "00", "00", "11", "00", "01", "11", "00", "11", "01", "01", "00", "00", "01", "01", "00", "11", "11", "01", "11", "00", "11", "01"),
302 => ("00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "00", "01", "11", "01", "00", "01", "11", "01", "11", "01", "11", "00", "11", "01", "00", "00", "01", "01", "00", "11", "00", "01"),
303 => ("01", "00", "00", "01", "00", "11", "11", "00", "00", "01", "11", "01", "11", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "00", "00", "01", "00"),
304 => ("00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "01", "00", "01", "11", "00", "00", "01", "00", "01", "01", "01", "01", "00", "11", "00", "11", "01", "00", "11", "11", "11"),
305 => ("00", "00", "01", "00", "00", "11", "11", "00", "01", "01", "00", "01", "00", "11", "00", "11", "01", "01", "01", "00", "11", "01", "01", "00", "01", "00", "11", "00", "01", "11", "01", "01"),
306 => ("01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "11", "11", "01", "01", "00", "00", "11", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "11"),
307 => ("00", "01", "00", "11", "00", "01", "01", "11", "11", "01", "01", "00", "11", "11", "00", "00", "01", "01", "01", "01", "01", "11", "11", "00", "00", "00", "01", "01", "01", "01", "01", "00"),
308 => ("00", "00", "01", "11", "11", "00", "11", "00", "11", "01", "00", "01", "01", "00", "01", "01", "11", "11", "00", "00", "01", "00", "11", "00", "01", "01", "00", "11", "01", "00", "00", "00"),
309 => ("01", "11", "01", "01", "11", "01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01", "11", "01", "11", "11", "01", "01", "01", "00", "00", "01"),
310 => ("00", "00", "00", "01", "11", "00", "01", "00", "11", "00", "00", "00", "11", "00", "00", "00", "01", "11", "00", "00", "11", "01", "01", "11", "00", "01", "11", "01", "00", "01", "00", "01"),
311 => ("01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "11", "11", "01", "01", "01", "01", "00", "01", "01", "00", "01"),
312 => ("00", "11", "01", "00", "11", "00", "01", "00", "00", "11", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "00", "00", "00", "01", "01", "11", "01", "11", "00", "11", "00", "01"),
313 => ("00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "11", "01", "11", "01", "01", "00", "11", "11", "00"),
314 => ("00", "11", "01", "01", "00", "11", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "00", "11", "01", "11", "01", "01", "01", "11", "11", "01", "01", "00", "11", "00", "00", "00"),
315 => ("01", "01", "11", "00", "11", "00", "11", "01", "11", "00", "00", "00", "01", "11", "11", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "00"),
316 => ("00", "01", "01", "00", "11", "00", "11", "01", "00", "01", "01", "00", "01", "01", "00", "01", "11", "11", "01", "01", "01", "01", "11", "01", "11", "00", "00", "11", "00", "00", "11", "01"),
317 => ("00", "11", "00", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "00", "11", "11", "00", "11", "00", "00", "01", "00", "01", "11", "00", "00", "00", "11", "00"),
318 => ("01", "11", "00", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "11", "11", "01", "00", "11", "00", "11", "00", "01", "00", "11", "01", "01"),
319 => ("01", "01", "01", "11", "00", "01", "11", "00", "11", "00", "00", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "11", "00", "00", "00", "11", "11", "00"),
320 => ("00", "00", "11", "01", "11", "01", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00", "11", "00", "01", "00", "11", "11", "01", "01", "00", "01", "00", "00", "11", "11", "01", "00"),
321 => ("01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "11", "01", "00", "01", "01", "00", "01", "11", "11", "01", "00", "00", "01", "01", "11", "01", "01", "11"),
322 => ("01", "00", "11", "01", "01", "00", "11", "00", "11", "01", "11", "01", "00", "00", "01", "01", "00", "00", "00", "11", "11", "01", "01", "11", "00", "01", "00", "11", "00", "00", "00", "00"),
323 => ("01", "11", "00", "11", "01", "00", "00", "00", "01", "11", "11", "01", "01", "00", "01", "00", "01", "11", "11", "01", "01", "01", "01", "01", "00", "01", "01", "00", "00", "11", "01", "11"),
324 => ("00", "11", "01", "00", "11", "00", "01", "01", "11", "11", "11", "01", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "00", "01", "00", "00", "01", "00", "00", "11"),
325 => ("00", "00", "01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "11", "11", "01", "11", "01", "11", "11", "01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "01"),
326 => ("01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "00", "01", "11", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "01", "11", "01", "01", "11", "00", "01", "00"),
327 => ("00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "11", "11", "00", "01", "00", "11", "11", "11", "01", "01", "01", "00", "00", "11", "00", "11", "00"),
328 => ("01", "01", "00", "01", "11", "01", "00", "00", "00", "11", "01", "11", "01", "01", "01", "00", "11", "00", "11", "01", "00", "11", "01", "00", "00", "00", "00", "01", "01", "11", "00", "11"),
329 => ("00", "00", "11", "01", "11", "11", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "11", "00", "00"),
330 => ("00", "01", "11", "00", "00", "01", "00", "11", "00", "01", "01", "01", "01", "00", "11", "01", "11", "00", "00", "00", "01", "11", "01", "01", "11", "00", "00", "00", "01", "01", "11", "11"),
331 => ("00", "00", "00", "01", "00", "00", "11", "11", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "01", "00", "00", "11", "11", "11", "00", "00", "01", "01", "01", "01", "11"),
332 => ("01", "11", "00", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "11", "00", "11", "00", "00", "00", "01", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00"),
333 => ("01", "00", "11", "00", "01", "00", "00", "00", "01", "11", "00", "00", "00", "01", "11", "00", "00", "01", "00", "11", "01", "11", "11", "11", "00", "00", "00", "00", "01", "00", "00", "00"),
334 => ("01", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "11", "01", "11", "00", "01", "11", "11", "11", "01", "00", "01", "11", "00", "00", "00", "00"),
335 => ("00", "01", "11", "00", "00", "01", "11", "00", "00", "00", "01", "11", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "00"),
336 => ("01", "01", "01", "01", "11", "01", "11", "11", "01", "00", "00", "00", "11", "11", "00", "00", "01", "00", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "00", "11", "01"),
337 => ("00", "11", "11", "01", "11", "01", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "11", "11", "11", "00"),
338 => ("01", "11", "00", "00", "01", "11", "11", "01", "00", "00", "00", "01", "01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "01", "11", "11", "01", "11", "00", "00", "00", "01", "00"),
339 => ("00", "01", "00", "11", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00", "11", "00", "01", "11", "00", "00", "11", "01", "01", "01", "01", "00", "01", "00", "00", "00"),
340 => ("00", "11", "01", "01", "11", "01", "01", "11", "01", "00", "11", "00", "00", "00", "00", "01", "01", "01", "01", "01", "11", "01", "00", "11", "00", "11", "11", "00", "00", "00", "00", "00"),
341 => ("01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "00", "11", "01", "11", "01", "01", "11", "00", "11", "00", "00", "01", "00", "11", "01", "11", "00", "01", "00", "00", "00"),
342 => ("01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "11", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "01", "11", "00", "01", "11", "01"),
343 => ("00", "00", "01", "01", "01", "11", "11", "00", "00", "00", "11", "11", "11", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "11", "00", "01", "01"),
344 => ("00", "01", "00", "11", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00", "11", "01", "00", "11", "01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "00", "11", "00"),
345 => ("01", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "00", "11", "01", "00", "11", "01", "00", "01", "00", "00", "01", "11", "00"),
346 => ("00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "00", "11", "01", "11", "00", "00", "00", "01", "11", "01", "00", "01", "00", "11", "11", "01", "11", "00", "01", "01"),
347 => ("01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "11", "01", "00", "01", "01", "00", "11", "11", "11", "01", "00", "01", "01", "11", "11"),
348 => ("00", "00", "11", "11", "11", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00"),
349 => ("01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "00", "00", "11", "00", "00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "01", "01", "01", "00", "01", "00", "11", "11"),
350 => ("01", "01", "00", "01", "01", "11", "11", "01", "00", "01", "00", "11", "11", "11", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11"),
351 => ("00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "11", "11", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00"),
352 => ("00", "00", "01", "00", "01", "00", "11", "11", "11", "01", "00", "01", "00", "01", "01", "00", "00", "11", "11", "00", "11", "01", "00", "01", "01", "01", "00", "11", "00", "01", "01", "00"),
353 => ("00", "01", "01", "11", "01", "11", "01", "00", "11", "00", "01", "11", "01", "00", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00", "01", "01", "00", "11", "01", "11", "00"),
354 => ("00", "00", "01", "01", "00", "00", "01", "00", "00", "01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "00", "11", "01", "11", "11", "01", "00", "01", "00", "11", "01", "01", "01"),
355 => ("01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "11", "11", "01", "11", "00", "00", "11", "00", "00", "01", "00", "11", "00"),
356 => ("01", "00", "01", "01", "11", "11", "11", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "11", "01", "00", "01", "00", "00", "01", "00", "01", "00", "01", "11", "00"),
357 => ("01", "11", "00", "00", "00", "01", "11", "11", "00", "00", "00", "11", "11", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "11", "01", "01"),
358 => ("01", "11", "00", "00", "00", "01", "11", "00", "11", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00"),
359 => ("00", "11", "00", "01", "00", "00", "11", "11", "00", "01", "00", "00", "11", "00", "11", "01", "01", "11", "00", "11", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "01", "00"),
360 => ("00", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "01", "01", "11", "00", "11", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "00", "01"),
361 => ("01", "00", "00", "11", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "01", "00", "00", "00", "01", "11", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "01", "11"),
362 => ("00", "00", "01", "11", "01", "11", "01", "01", "00", "11", "01", "00", "01", "11", "00", "01", "11", "00", "11", "00", "00", "01", "11", "11", "01", "01", "00", "00", "00", "00", "01", "01"),
363 => ("01", "00", "00", "00", "01", "11", "00", "11", "01", "11", "00", "11", "01", "00", "01", "00", "11", "00", "00", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "11", "00", "01"),
364 => ("00", "11", "01", "00", "11", "11", "11", "00", "11", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "00", "01", "01"),
365 => ("00", "00", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "11", "01", "01", "11", "01", "11", "01", "11", "00", "01", "00", "00", "11", "11", "01", "01", "00", "11"),
366 => ("00", "01", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "01", "00", "11", "00", "11", "01", "01", "00", "11", "00", "01", "11", "11", "00", "00", "00", "00", "11", "00"),
367 => ("01", "01", "01", "00", "00", "11", "00", "11", "01", "01", "11", "01", "11", "01", "00", "00", "01", "11", "00", "01", "11", "00", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01"),
368 => ("01", "11", "01", "01", "00", "11", "01", "01", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "11", "00", "01", "00", "00", "00", "01", "00", "01", "11", "11", "00", "11", "01"),
369 => ("00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "11", "01", "11", "00", "00", "11", "11", "01", "01", "01", "01", "00"),
370 => ("00", "01", "00", "00", "11", "00", "01", "11", "11", "01", "00", "00", "00", "11", "00", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11", "01", "00", "01", "01"),
371 => ("00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "00", "11", "01", "01", "00", "01", "11", "01", "01", "00", "11", "11", "11", "01", "11", "11", "01", "00", "00", "00", "00", "01"),
372 => ("00", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "01", "11", "01", "00", "00", "11", "11", "11", "01", "11", "00", "00", "01", "00", "00", "01", "00"),
373 => ("01", "11", "11", "01", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "00", "00", "01", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00", "00", "00"),
374 => ("01", "00", "00", "11", "01", "01", "00", "01", "00", "11", "00", "01", "11", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "01", "00", "11", "11"),
375 => ("00", "00", "11", "01", "00", "00", "00", "01", "11", "01", "01", "11", "01", "01", "00", "11", "01", "11", "11", "01", "11", "01", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00"),
376 => ("01", "00", "11", "00", "00", "11", "00", "00", "00", "11", "11", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "11", "00"),
377 => ("01", "00", "11", "11", "01", "11", "00", "11", "01", "00", "00", "11", "00", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "01", "01", "01"),
378 => ("00", "11", "00", "11", "01", "01", "11", "00", "00", "00", "00", "11", "11", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "11", "01", "00", "01"),
379 => ("01", "00", "01", "00", "11", "11", "00", "11", "00", "01", "01", "11", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "00", "01", "11", "00", "11", "00", "11", "01", "01", "01"),
380 => ("00", "01", "01", "11", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "01", "11", "01", "01", "11", "11", "11", "01", "01", "11", "01", "00", "01"),
381 => ("00", "01", "11", "01", "00", "01", "11", "11", "00", "00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "00", "11", "00", "11", "01", "00", "01", "00", "00", "01", "01"),
382 => ("01", "00", "11", "00", "11", "00", "11", "01", "11", "11", "00", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00", "00", "11", "00", "01", "01", "00"),
383 => ("01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "11", "00", "00", "00", "11", "01", "11", "11", "01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "00"),
384 => ("00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "11", "00", "01", "01", "01", "01", "00", "11", "01", "00", "11", "11", "11", "00", "00", "11", "00", "00", "00", "00", "00", "00"),
385 => ("00", "00", "11", "01", "01", "00", "11", "00", "01", "00", "00", "11", "01", "01", "00", "01", "00", "11", "00", "01", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01"),
386 => ("00", "11", "00", "11", "00", "11", "01", "01", "11", "00", "00", "01", "00", "01", "01", "01", "11", "00", "11", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "00"),
387 => ("00", "11", "01", "11", "00", "01", "00", "00", "11", "00", "00", "01", "11", "00", "01", "01", "00", "00", "11", "00", "11", "11", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00"),
388 => ("00", "00", "01", "01", "01", "11", "00", "00", "11", "01", "00", "11", "01", "01", "11", "01", "00", "01", "01", "00", "00", "00", "00", "11", "11", "11", "01", "01", "01", "01", "00", "00"),
389 => ("00", "01", "01", "01", "00", "11", "00", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "01", "11", "11", "01", "00", "01", "00", "11", "00", "01", "00", "11", "11", "00", "00"),
390 => ("00", "00", "11", "01", "00", "11", "11", "00", "01", "11", "00", "00", "01", "00", "11", "01", "11", "00", "00", "01", "11", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01"),
391 => ("01", "00", "00", "00", "01", "11", "11", "01", "11", "01", "01", "00", "00", "00", "01", "01", "11", "00", "01", "11", "00", "01", "01", "11", "01", "00", "01", "01", "00", "11", "11", "00"),
392 => ("01", "00", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "00", "11", "11", "00", "01", "01", "00", "11", "01", "00", "01", "11", "01", "01", "00", "01", "01", "01", "01"),
393 => ("00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "11", "00", "00", "11", "00", "11", "01", "01", "00", "11", "01", "00", "01", "11", "00", "11", "00", "01", "11", "00", "01", "00"),
394 => ("00", "01", "11", "01", "01", "11", "01", "11", "00", "01", "01", "11", "11", "00", "01", "11", "00", "01", "01", "11", "01", "01", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01"),
395 => ("00", "11", "11", "00", "00", "11", "01", "01", "00", "11", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11", "01", "01", "00", "00", "00", "01", "01", "11", "11", "11", "00"),
396 => ("01", "00", "00", "00", "01", "00", "11", "01", "00", "11", "11", "01", "00", "11", "00", "00", "00", "11", "01", "11", "00", "11", "01", "01", "11", "00", "00", "01", "00", "01", "01", "00"),
397 => ("01", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "11", "01", "00", "11", "00", "00", "01", "01", "00", "00", "00", "01", "01", "01", "00", "11", "01", "11"),
398 => ("00", "01", "01", "01", "00", "01", "00", "11", "11", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "01", "11", "11", "00", "01", "01", "00", "11", "00", "01", "01", "01", "00"),
399 => ("00", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "11", "11", "00", "00", "11", "00", "00", "00", "11", "00", "11", "01", "00", "00", "11", "01", "01", "00", "01", "00"),
400 => ("00", "00", "01", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "11", "11", "01", "00", "00", "01", "11", "00", "01", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01"),
401 => ("00", "11", "11", "11", "01", "01", "11", "00", "01", "01", "11", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01", "01", "00", "11", "01", "00", "11"),
402 => ("01", "11", "11", "01", "00", "01", "01", "00", "00", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "11", "00", "01", "01", "11", "01", "11"),
403 => ("01", "01", "00", "00", "00", "01", "11", "00", "01", "11", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "11", "11", "01", "00", "01", "01", "00", "11", "01", "01"),
404 => ("01", "01", "11", "01", "11", "00", "11", "01", "01", "11", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "00"),
405 => ("00", "11", "01", "00", "00", "11", "01", "11", "00", "01", "11", "00", "11", "01", "01", "00", "01", "00", "01", "00", "11", "11", "00", "11", "01", "01", "01", "00", "00", "00", "00", "01"),
406 => ("01", "01", "11", "00", "01", "01", "00", "11", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "11", "00", "00", "11", "00", "00", "11", "01", "00", "11"),
407 => ("00", "01", "11", "00", "01", "00", "11", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "11"),
408 => ("01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "11", "00", "00", "01", "11", "00", "00", "01", "01", "01", "00", "11", "00", "11", "00", "11", "01", "00", "11"),
409 => ("00", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "11", "00", "00", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "00", "11", "00", "01", "11"),
410 => ("00", "01", "00", "01", "00", "00", "11", "01", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "00", "11", "00", "11", "01", "11", "01", "01"),
411 => ("00", "11", "01", "00", "01", "00", "01", "01", "00", "11", "11", "01", "01", "01", "11", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "11", "11", "11"),
412 => ("00", "00", "01", "00", "01", "00", "00", "00", "11", "11", "11", "00", "01", "11", "00", "01", "11", "01", "11", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "01", "00"),
413 => ("01", "01", "01", "00", "00", "00", "11", "11", "00", "11", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "00", "00", "11", "11"),
414 => ("00", "11", "00", "11", "01", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "11", "11", "00", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "01", "01", "00", "11"),
415 => ("00", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "11", "00", "11", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01"),
416 => ("01", "01", "01", "01", "01", "00", "01", "11", "11", "00", "11", "01", "00", "01", "11", "01", "01", "11", "00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01"),
417 => ("01", "01", "01", "01", "00", "01", "11", "01", "01", "00", "11", "00", "11", "01", "01", "00", "11", "00", "00", "11", "01", "11", "01", "01", "11", "01", "01", "01", "11", "00", "00", "01"),
418 => ("01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "11", "00", "11", "01", "01", "11", "00", "00", "00", "00", "00", "01", "11", "01", "11", "01", "11", "00", "00", "00", "00", "00"),
419 => ("00", "01", "11", "01", "01", "01", "01", "01", "11", "11", "01", "01", "01", "00", "00", "00", "00", "01", "01", "11", "01", "01", "11", "01", "01", "01", "11", "11", "00", "00", "01", "01"),
420 => ("00", "00", "01", "00", "00", "11", "01", "00", "11", "01", "11", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "01", "11", "01", "01", "11", "01", "00"),
421 => ("00", "01", "11", "00", "01", "00", "01", "01", "00", "01", "00", "01", "00", "11", "11", "11", "11", "01", "00", "11", "00", "01", "11", "01", "00", "00", "01", "01", "11", "01", "00", "01"),
422 => ("00", "01", "01", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "11", "01", "00", "01", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00", "11"),
423 => ("00", "01", "00", "11", "01", "11", "00", "11", "00", "00", "01", "00", "01", "00", "01", "00", "01", "11", "00", "01", "00", "00", "11", "01", "11", "00", "00", "00", "01", "01", "01", "01"),
424 => ("00", "11", "11", "11", "01", "00", "00", "01", "00", "01", "11", "11", "01", "00", "00", "11", "00", "00", "11", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "01", "01"),
425 => ("00", "01", "01", "01", "00", "00", "00", "11", "11", "00", "00", "11", "11", "01", "00", "01", "01", "01", "11", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "11", "00"),
426 => ("00", "00", "01", "00", "01", "11", "00", "00", "11", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "11", "00", "00", "00", "11"),
427 => ("01", "11", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "11", "11", "01", "01", "11", "01", "11", "00", "00", "00", "11", "11", "00", "01"),
428 => ("01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "11", "00", "00", "00", "01", "00", "00", "11", "01", "11", "00", "01", "11", "01", "00", "01", "00", "11", "01", "00", "00", "11"),
429 => ("00", "11", "01", "11", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "00", "11", "01", "00", "11", "00"),
430 => ("01", "00", "00", "00", "00", "01", "11", "00", "00", "11", "01", "11", "00", "11", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "00"),
431 => ("01", "11", "00", "11", "00", "01", "00", "11", "00", "01", "11", "01", "00", "00", "00", "00", "01", "11", "00", "11", "01", "01", "00", "00", "00", "01", "01", "00", "01", "01", "11", "00"),
432 => ("01", "00", "00", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "00", "11", "01", "11", "01", "11", "11", "01", "00", "00", "01", "11", "01", "00"),
433 => ("01", "11", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "01", "00", "00", "11", "01", "00", "11", "11", "01", "01", "01", "11", "01", "01"),
434 => ("00", "01", "00", "00", "01", "11", "01", "11", "11", "00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "01", "11", "00"),
435 => ("01", "01", "11", "00", "00", "01", "01", "11", "11", "01", "01", "00", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "00", "01", "01", "01", "01", "11", "00", "00"),
436 => ("00", "11", "01", "11", "11", "00", "00", "01", "00", "01", "01", "00", "11", "01", "01", "01", "11", "11", "00", "00", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "11", "01"),
437 => ("00", "01", "01", "01", "00", "00", "11", "01", "11", "00", "11", "01", "01", "11", "00", "01", "01", "11", "11", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "01", "01", "01"),
438 => ("01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "11", "11", "11", "11", "11", "01", "01", "00", "00", "00", "01", "00", "00", "00"),
439 => ("00", "00", "01", "11", "11", "11", "01", "01", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00"),
440 => ("00", "00", "01", "11", "11", "00", "11", "01", "11", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "00", "00"),
441 => ("01", "11", "00", "01", "11", "01", "01", "01", "11", "00", "01", "00", "11", "00", "11", "00", "00", "01", "00", "00", "01", "00", "00", "01", "00", "01", "11", "00", "11", "00", "01", "01"),
442 => ("01", "11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "00", "11", "11", "01", "01"),
443 => ("01", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "00", "00", "11", "01", "01", "11", "01", "01", "11", "00", "11", "00", "11", "01", "01", "11", "00", "01", "00", "11", "01"),
444 => ("01", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "00", "11", "00", "01", "00", "11", "01", "01", "11", "00", "11", "00", "01", "11", "00", "11", "00", "11", "01", "01"),
445 => ("01", "01", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "11", "11", "11", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "11", "01", "00", "00", "00", "00", "11"),
446 => ("01", "00", "00", "00", "00", "00", "11", "00", "00", "11", "11", "01", "11", "00", "01", "11", "00", "11", "00", "11", "00", "01", "01", "11", "01", "01", "00", "00", "00", "00", "00", "00"),
447 => ("00", "00", "01", "11", "00", "11", "01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "01", "11", "01", "01", "11", "01", "01", "11", "00", "01", "01", "01", "01", "11", "01"),
448 => ("01", "11", "01", "01", "00", "00", "11", "11", "00", "00", "00", "11", "11", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "11", "11", "01", "00", "00", "01", "01", "01", "01"),
449 => ("01", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "01", "11", "01", "00", "01", "00", "01", "00", "11", "11", "00", "00", "01", "00", "11", "00", "01", "01", "11", "11", "01"),
450 => ("01", "00", "01", "11", "01", "11", "01", "00", "11", "01", "11", "01", "01", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "01", "11", "00", "01"),
451 => ("01", "11", "11", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "11", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "11", "00", "01", "11"),
452 => ("00", "00", "11", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "11", "01", "01", "00", "11", "01", "01", "11", "00", "00", "11", "01", "01", "00", "01", "01", "00"),
453 => ("01", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "00", "00", "01", "11", "11", "11", "11", "01", "00", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "00", "11"),
454 => ("01", "01", "01", "00", "11", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "11", "01", "11", "01", "00", "11", "01", "01", "11", "00"),
455 => ("00", "01", "01", "01", "01", "00", "01", "11", "11", "01", "11", "11", "01", "11", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "11", "01", "00"),
456 => ("01", "00", "11", "00", "01", "11", "11", "00", "01", "00", "11", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "00", "01", "00", "11", "00", "00", "11", "01", "00", "01"),
457 => ("01", "11", "00", "01", "00", "01", "11", "11", "11", "11", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "00", "00", "11", "01", "01", "01", "00", "11", "00", "00"),
458 => ("01", "00", "00", "11", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "00", "00", "11", "00", "11", "00", "11", "00", "01", "11", "01", "01", "00", "00"),
459 => ("00", "11", "01", "01", "11", "11", "01", "11", "01", "11", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "01", "00", "11", "11", "01", "01", "01", "00"),
460 => ("00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "00", "01", "00", "11", "00", "11", "11", "00", "00", "11", "11", "00", "00", "00", "01", "00", "01", "11", "01", "01"),
461 => ("00", "01", "11", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "00", "11", "01", "01", "01", "01", "11", "01", "00", "11"),
462 => ("00", "00", "01", "01", "01", "11", "11", "00", "01", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "11", "01", "00"),
463 => ("00", "01", "01", "01", "01", "11", "00", "01", "00", "11", "00", "11", "11", "01", "00", "11", "11", "11", "00", "01", "00", "00", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
464 => ("00", "01", "11", "00", "00", "11", "00", "00", "00", "11", "01", "01", "00", "00", "00", "11", "00", "11", "11", "00", "11", "01", "00", "00", "00", "01", "01", "11", "01", "01", "01", "00"),
465 => ("01", "00", "01", "00", "11", "01", "01", "00", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "11", "01", "11", "01", "11", "01", "00", "00", "11", "11", "00"),
466 => ("01", "01", "01", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "11", "00", "01", "00", "11", "00", "01", "01", "11", "11", "01", "01", "11", "01", "00"),
467 => ("01", "11", "00", "01", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "11", "00", "00", "11", "01", "00", "00"),
468 => ("01", "00", "01", "00", "00", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "11", "01", "00", "00", "00", "00", "11", "01", "01", "11", "00", "11", "00", "11", "01", "01", "11"),
469 => ("00", "01", "01", "01", "00", "01", "01", "00", "11", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "00", "11", "00", "00", "01", "11", "11", "01", "01", "11", "00"),
470 => ("01", "11", "11", "01", "01", "01", "11", "01", "11", "01", "00", "01", "01", "11", "11", "01", "01", "00", "01", "01", "01", "01", "00", "01", "01", "00", "01", "11", "11", "01", "00", "01"),
471 => ("00", "00", "00", "01", "00", "01", "00", "01", "00", "01", "00", "11", "00", "11", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "11", "01", "11", "00", "00", "00", "11", "00"),
472 => ("00", "11", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", "01", "11", "00", "00", "00", "01", "01", "00", "11", "01"),
473 => ("00", "01", "00", "11", "01", "00", "01", "11", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "11", "01", "00", "00", "11", "00", "11", "01", "11", "01", "01"),
474 => ("00", "01", "01", "00", "01", "00", "11", "01", "01", "01", "00", "11", "01", "01", "00", "11", "01", "11", "01", "00", "00", "11", "01", "01", "11", "11", "01", "01", "00", "00", "00", "01"),
475 => ("00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "11", "00", "11", "11", "01", "00", "00", "01", "00", "01", "11", "00", "00", "00", "00"),
476 => ("01", "11", "11", "01", "00", "01", "11", "11", "11", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "00", "11", "11", "01", "01", "00", "01", "00", "01", "00", "00", "00", "00"),
477 => ("00", "00", "01", "11", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "01", "01", "11", "11", "01", "01", "00", "01", "11", "11", "00"),
478 => ("01", "11", "01", "00", "00", "00", "11", "11", "00", "01", "11", "11", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "11", "01", "01", "00", "01"),
479 => ("00", "01", "00", "01", "00", "01", "01", "11", "11", "00", "01", "11", "00", "11", "00", "00", "00", "00", "11", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "00", "00", "11"),
480 => ("00", "00", "11", "01", "11", "00", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "11", "11", "11"),
481 => ("00", "00", "00", "01", "11", "11", "01", "01", "11", "11", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "00", "11", "01", "00", "00", "11", "00", "01", "01", "01", "01", "00"),
482 => ("01", "01", "11", "00", "00", "00", "00", "01", "00", "11", "01", "00", "00", "01", "00", "11", "00", "00", "11", "11", "01", "00", "11", "01", "11", "00", "00", "00", "11", "00", "01", "01"),
483 => ("01", "11", "00", "00", "01", "00", "01", "01", "00", "11", "11", "00", "01", "11", "00", "11", "01", "00", "01", "01", "11", "00", "11", "01", "00", "01", "01", "00", "00", "11", "00", "01"),
484 => ("00", "11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "00", "01", "01", "00", "00", "11", "11", "11", "00", "01", "00", "00", "11", "01", "11", "00", "11", "01", "01", "01"),
485 => ("01", "01", "11", "11", "11", "01", "00", "00", "11", "01", "11", "01", "00", "01", "11", "01", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "11", "01", "00", "00"),
486 => ("01", "11", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "11", "01", "01", "11", "01", "00", "11", "00", "00", "00", "11", "01", "11", "01", "00"),
487 => ("01", "00", "01", "01", "01", "11", "01", "00", "11", "11", "00", "00", "01", "00", "11", "11", "00", "01", "01", "11", "00", "01", "00", "00", "11", "00", "11", "00", "00", "00", "00", "01"),
488 => ("01", "11", "00", "00", "00", "00", "11", "01", "11", "01", "00", "00", "00", "01", "00", "01", "01", "00", "01", "11", "11", "00", "01", "01", "00", "01", "01", "11", "00", "11", "01", "00"),
489 => ("01", "01", "01", "00", "01", "01", "11", "01", "11", "00", "00", "01", "11", "01", "11", "01", "00", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "00", "00", "00", "00", "11"),
490 => ("01", "00", "01", "01", "01", "00", "01", "11", "00", "11", "00", "01", "01", "01", "00", "11", "11", "00", "01", "00", "11", "00", "01", "11", "01", "00", "11", "00", "01", "00", "00", "01"),
491 => ("01", "01", "11", "00", "01", "11", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01"),
492 => ("01", "00", "01", "11", "01", "00", "01", "00", "01", "00", "00", "00", "01", "00", "11", "11", "00", "01", "00", "01", "01", "01", "01", "11", "01", "11", "00", "11", "00", "01", "01", "11"),
493 => ("00", "00", "11", "00", "01", "11", "00", "01", "11", "01", "01", "11", "11", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "11", "00"),
494 => ("01", "00", "01", "11", "01", "01", "01", "00", "11", "00", "11", "11", "11", "00", "00", "00", "00", "11", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "01", "01", "00"),
495 => ("01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "11", "11", "00", "11", "00", "01", "00", "11", "01", "11", "01", "11", "01", "01", "01", "11", "11", "01", "01"),
496 => ("00", "11", "01", "00", "01", "00", "11", "01", "11", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "11", "01", "00", "01", "11", "01", "01", "01", "00", "01", "01", "01"),
497 => ("01", "00", "00", "01", "11", "01", "00", "00", "00", "00", "11", "01", "11", "00", "01", "01", "00", "11", "01", "00", "11", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01"),
498 => ("00", "01", "00", "01", "00", "11", "00", "11", "11", "01", "00", "01", "11", "01", "00", "00", "01", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01", "11", "11", "00", "01", "00"),
499 => ("00", "11", "01", "00", "01", "01", "00", "01", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "11", "00", "00", "00", "00", "11", "01", "01", "11", "01", "01", "01", "01", "11")),
(
0 => ("01", "00", "01", "01", "00", "00", "01", "11", "01", "11", "00", "11", "01", "00", "00", "01", "11", "01", "01", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "11", "00", "01"),
1 => ("00", "00", "00", "01", "00", "01", "00", "00", "11", "01", "11", "01", "11", "01", "01", "00", "11", "01", "01", "00", "01", "11", "01", "00", "11", "01", "11", "11", "01", "01", "01", "01"),
2 => ("00", "11", "11", "01", "11", "01", "11", "11", "00", "11", "01", "01", "01", "01", "01", "11", "01", "00", "01", "00", "11", "01", "01", "00", "01", "00", "00", "01", "01", "00", "00", "11"),
3 => ("00", "01", "00", "01", "11", "11", "01", "01", "11", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "00", "11", "00", "01", "00", "01", "11", "01", "01"),
4 => ("01", "01", "11", "01", "11", "11", "01", "00", "00", "11", "01", "11", "00", "00", "11", "11", "01", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "00", "11", "00", "00"),
5 => ("01", "00", "11", "01", "01", "01", "00", "00", "00", "11", "00", "01", "01", "00", "11", "00", "01", "11", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "11", "11", "01"),
6 => ("01", "11", "11", "11", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "00", "00", "11", "00", "01", "11", "00", "11", "00", "01", "01", "00", "00", "11", "11", "00", "01", "00"),
7 => ("01", "11", "00", "11", "00", "01", "01", "01", "11", "01", "11", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "00", "11", "01", "11", "00", "00", "11", "01", "01", "01", "11"),
8 => ("00", "11", "11", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "00", "00", "00", "11", "11", "01", "01", "11", "01", "01", "01", "01", "11", "11", "00"),
9 => ("00", "11", "01", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "01", "01", "01", "11", "00", "11", "01", "11", "01", "01", "01", "01", "11", "00", "01", "01", "11", "01"),
10 => ("01", "01", "00", "00", "01", "01", "00", "11", "01", "01", "00", "11", "11", "00", "00", "01", "11", "00", "01", "01", "11", "01", "11", "00", "01", "00", "00", "01", "11", "11", "01", "01"),
11 => ("00", "01", "00", "11", "11", "11", "00", "11", "01", "00", "11", "00", "00", "00", "01", "01", "11", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01"),
12 => ("00", "00", "00", "00", "00", "01", "01", "11", "00", "11", "00", "01", "11", "11", "00", "01", "01", "01", "00", "11", "01", "01", "11", "00", "00", "00", "01", "00", "00", "00", "11", "01"),
13 => ("00", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "11", "00", "11", "11", "11", "01", "00", "00", "00", "01", "11", "11", "00", "01", "01", "00", "00", "00", "01", "00", "11"),
14 => ("01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "00", "11", "01", "01", "01", "11", "11", "00", "11", "00", "11", "11", "00"),
15 => ("00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "11", "00", "00", "01", "11", "00", "11", "11", "11", "11", "01", "00", "00", "00", "01", "01", "00", "11", "01", "00", "11", "00"),
16 => ("01", "01", "00", "01", "01", "11", "00", "01", "00", "01", "11", "00", "01", "01", "11", "01", "01", "11", "00", "00", "01", "11", "00", "01", "01", "00", "01", "11", "00", "01", "11", "01"),
17 => ("01", "11", "11", "11", "00", "11", "00", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "11", "00", "00", "01", "00", "00", "01", "00", "00", "11", "01", "01", "00"),
18 => ("01", "11", "01", "00", "01", "11", "00", "01", "00", "00", "01", "01", "11", "01", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "11", "11", "11", "01", "01", "01"),
19 => ("00", "01", "01", "11", "11", "01", "01", "01", "11", "01", "00", "11", "00", "01", "01", "11", "01", "01", "01", "00", "01", "11", "01", "00", "01", "00", "11", "11", "00", "00", "00", "01"),
20 => ("01", "00", "01", "01", "00", "01", "11", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "01", "00", "11", "00", "11", "00", "11"),
21 => ("00", "11", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "11", "00", "00", "11", "11", "00", "00", "00", "01", "11", "11", "01", "00", "01", "00", "11"),
22 => ("01", "01", "11", "00", "11", "00", "01", "01", "00", "01", "00", "00", "11", "01", "01", "01", "00", "00", "00", "01", "01", "11", "11", "01", "01", "01", "01", "11", "00", "00", "11", "11"),
23 => ("00", "00", "11", "00", "00", "00", "01", "11", "00", "01", "00", "01", "11", "01", "00", "00", "00", "01", "00", "11", "11", "01", "00", "11", "11", "00", "00", "01", "01", "11", "00", "11"),
24 => ("00", "01", "00", "11", "00", "00", "00", "01", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "01", "11", "00", "01", "01", "11", "01", "00", "01", "11", "00", "11", "00", "11"),
25 => ("01", "11", "00", "11", "01", "01", "11", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "00", "00", "01", "11", "11", "00", "00", "11", "00"),
26 => ("01", "01", "00", "11", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "11", "11", "00", "11", "01", "00", "11", "01", "11", "11"),
27 => ("00", "00", "01", "11", "01", "11", "11", "00", "01", "01", "00", "00", "00", "11", "00", "00", "01", "11", "00", "00", "00", "01", "01", "00", "11", "01", "11", "11", "00", "01", "00", "00"),
28 => ("00", "01", "00", "01", "11", "01", "01", "00", "01", "11", "01", "11", "00", "00", "00", "01", "00", "01", "11", "00", "00", "01", "01", "11", "11", "00", "11", "01", "00", "01", "00", "01"),
29 => ("00", "01", "01", "01", "01", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "01", "11", "01", "01", "11", "01", "00", "11", "01", "00", "11", "11", "01", "01", "01", "01", "11"),
30 => ("00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "00", "00", "11", "01", "00", "01", "00", "01", "00", "11", "11", "11", "00", "00", "00", "11", "01", "11", "11", "00", "01", "00"),
31 => ("00", "01", "00", "11", "01", "01", "11", "00", "00", "11", "01", "00", "00", "00", "11", "00", "01", "00", "11", "01", "00", "11", "00", "00", "01", "01", "11", "11", "01", "01", "01", "00"),
32 => ("01", "11", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "00", "11", "00", "11", "01", "11", "00", "11", "00", "11", "01", "00", "11", "00", "00", "11", "01", "00", "01", "11"),
33 => ("00", "00", "01", "11", "11", "00", "01", "01", "01", "11", "01", "01", "00", "00", "11", "11", "01", "00", "00", "01", "11", "11", "11", "00", "01", "00", "11", "01", "01", "01", "01", "01"),
34 => ("01", "11", "11", "11", "11", "01", "01", "01", "00", "00", "00", "01", "11", "00", "00", "00", "11", "00", "00", "00", "11", "11", "01", "01", "00", "00", "00", "00", "11", "01", "00", "00"),
35 => ("00", "11", "00", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "01", "00", "11", "01", "11", "00", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "11", "11", "00"),
36 => ("00", "01", "00", "01", "01", "00", "00", "11", "11", "00", "01", "11", "11", "11", "01", "11", "11", "01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "01", "01", "00", "00", "11"),
37 => ("01", "01", "11", "00", "00", "01", "01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "00", "11", "11", "00", "01", "00", "01", "00", "11", "01", "11", "01", "00", "00", "11", "11"),
38 => ("01", "01", "11", "01", "11", "00", "00", "00", "11", "00", "01", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "11", "00", "00", "11", "01", "01", "00", "11", "01", "00", "00"),
39 => ("01", "01", "11", "00", "11", "01", "11", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "00", "11", "00", "00", "00", "01", "00", "01", "11", "11", "01", "01"),
40 => ("01", "11", "11", "01", "00", "11", "01", "00", "11", "01", "11", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "11", "00", "11", "00", "00", "01", "00", "01", "11", "01", "01"),
41 => ("01", "01", "00", "00", "01", "00", "01", "11", "01", "00", "11", "01", "11", "00", "01", "00", "01", "01", "11", "00", "01", "11", "01", "11", "00", "11", "01", "00", "01", "00", "11", "01"),
42 => ("00", "11", "11", "01", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "01"),
43 => ("01", "01", "01", "11", "00", "11", "00", "11", "01", "00", "11", "00", "00", "01", "11", "01", "11", "01", "00", "01", "00", "01", "00", "11", "00", "11", "00", "01", "00", "01", "11", "01"),
44 => ("01", "00", "00", "00", "11", "11", "11", "01", "00", "01", "11", "00", "00", "01", "00", "11", "01", "01", "00", "11", "01", "01", "00", "00", "00", "11", "01", "00", "00", "00", "00", "01"),
45 => ("00", "00", "11", "11", "11", "01", "01", "11", "11", "00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "11", "11", "01", "11", "00", "00", "01", "01", "01"),
46 => ("00", "01", "00", "11", "11", "00", "11", "00", "00", "00", "11", "11", "11", "00", "00", "01", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "00", "01", "00", "11", "01", "00"),
47 => ("01", "11", "01", "00", "11", "01", "01", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "00", "11", "01", "01", "00", "01", "11", "01", "01", "11", "01", "11", "11", "00", "01"),
48 => ("01", "00", "00", "01", "11", "11", "00", "11", "00", "11", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "11", "01", "00", "11", "00", "01", "01", "00", "11", "00", "01", "00"),
49 => ("00", "00", "11", "01", "01", "00", "01", "00", "01", "11", "11", "11", "00", "00", "01", "11", "00", "01", "01", "00", "00", "01", "00", "01", "01", "01", "01", "01", "00", "11", "00", "11"),
50 => ("00", "11", "01", "00", "01", "11", "00", "01", "00", "01", "00", "00", "00", "11", "00", "01", "00", "00", "00", "01", "00", "11", "01", "01", "11", "01", "11", "11", "01", "00", "01", "01"),
51 => ("00", "01", "01", "11", "01", "11", "00", "01", "01", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01", "00", "11", "01", "00", "00", "01", "00", "11", "00", "00", "01", "11", "11"),
52 => ("01", "11", "00", "00", "00", "00", "11", "00", "11", "11", "11", "00", "11", "00", "00", "01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00"),
53 => ("00", "01", "11", "11", "11", "00", "00", "01", "11", "00", "00", "00", "00", "11", "01", "11", "01", "11", "01", "00", "01", "11", "01", "00", "00", "00", "01", "11", "01", "00", "01", "00"),
54 => ("01", "01", "01", "01", "11", "01", "00", "01", "01", "11", "11", "00", "11", "00", "11", "00", "01", "11", "01", "00", "11", "01", "00", "00", "00", "00", "00", "01", "00", "00", "01", "11"),
55 => ("00", "00", "00", "00", "11", "01", "01", "00", "01", "01", "11", "11", "00", "00", "01", "01", "01", "01", "00", "11", "00", "00", "01", "01", "11", "11", "11", "01", "11", "01", "00", "01"),
56 => ("00", "00", "11", "11", "00", "11", "01", "11", "00", "11", "00", "00", "01", "00", "11", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "11", "01", "00"),
57 => ("00", "01", "01", "00", "01", "01", "01", "00", "01", "11", "01", "11", "00", "00", "00", "11", "00", "11", "01", "01", "01", "00", "00", "01", "00", "00", "11", "00", "00", "11", "11", "00"),
58 => ("01", "01", "01", "11", "01", "11", "00", "01", "01", "11", "01", "00", "11", "01", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "00", "11", "01", "11", "11", "01", "00", "00"),
59 => ("00", "01", "11", "11", "01", "00", "00", "01", "11", "01", "00", "11", "01", "01", "01", "11", "01", "11", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "11", "00", "00", "01"),
60 => ("00", "01", "01", "00", "11", "01", "00", "01", "00", "01", "00", "11", "01", "11", "01", "11", "01", "00", "00", "11", "01", "01", "00", "11", "01", "00", "11", "01", "01", "11", "00", "01"),
61 => ("01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "11", "11", "01", "01", "11", "01", "01", "00", "00", "11", "11", "01", "00", "00", "11", "11", "00", "11", "01", "00", "00", "00"),
62 => ("01", "11", "00", "01", "00", "00", "00", "00", "11", "11", "01", "00", "01", "11", "11", "00", "00", "01", "01", "01", "11", "11", "01", "00", "00", "00", "11", "00", "00", "11", "01", "00"),
63 => ("00", "00", "00", "01", "01", "00", "11", "11", "00", "00", "01", "11", "01", "00", "01", "00", "11", "00", "01", "01", "01", "11", "01", "00", "01", "11", "00", "01", "11", "11", "00", "11"),
64 => ("01", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "00", "11", "00", "11", "11", "11"),
65 => ("01", "01", "01", "00", "00", "01", "00", "00", "01", "11", "00", "11", "11", "01", "01", "00", "00", "01", "00", "11", "11", "00", "11", "00", "00", "11", "01", "11", "11", "00", "01", "00"),
66 => ("01", "00", "00", "01", "11", "00", "01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "01", "11", "11", "00", "01", "00", "00", "01", "11", "00", "11", "00", "00", "00", "00"),
67 => ("01", "00", "00", "01", "00", "00", "11", "11", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "11", "01", "00", "11", "11", "00", "01", "11", "00", "01", "11", "01", "00", "00"),
68 => ("01", "00", "00", "01", "00", "00", "11", "11", "00", "00", "01", "00", "00", "00", "01", "01", "01", "00", "00", "11", "11", "00", "11", "01", "00", "01", "00", "11", "11", "00", "11", "00"),
69 => ("00", "01", "11", "00", "01", "00", "01", "11", "11", "01", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "11", "11", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11"),
70 => ("01", "11", "11", "11", "00", "11", "11", "01", "11", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "01", "11", "01", "01", "01", "01", "01", "01", "01", "00", "01", "11", "01"),
71 => ("01", "11", "00", "00", "00", "01", "01", "01", "11", "11", "00", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "01", "01", "00"),
72 => ("01", "11", "01", "01", "00", "01", "11", "01", "00", "00", "00", "01", "11", "01", "11", "00", "00", "00", "11", "00", "01", "01", "11", "11", "11", "01", "00", "01", "01", "01", "01", "01"),
73 => ("01", "00", "01", "11", "00", "00", "11", "01", "01", "11", "00", "00", "11", "11", "11", "00", "00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "00", "01", "00", "01", "01", "00"),
74 => ("00", "01", "11", "01", "11", "01", "01", "00", "00", "01", "11", "00", "00", "00", "00", "00", "01", "01", "11", "00", "00", "00", "11", "00", "00", "11", "01", "11", "01", "01", "11", "01"),
75 => ("01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "11", "01", "00", "01", "01", "01", "00", "01", "00", "01", "11", "11", "00", "11", "11", "11", "01", "00", "01", "11", "01", "01"),
76 => ("00", "00", "01", "00", "00", "11", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "11", "01", "00", "11", "00", "11", "11", "00", "11", "11", "00", "00", "01", "01", "00", "11"),
77 => ("01", "00", "01", "00", "00", "11", "11", "00", "00", "01", "01", "11", "01", "01", "00", "01", "00", "11", "01", "11", "00", "00", "11", "11", "01", "00", "11", "01", "01", "01", "00", "00"),
78 => ("01", "11", "11", "00", "01", "01", "11", "11", "11", "11", "00", "01", "01", "01", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "00", "01", "11", "11", "00", "01", "00", "01"),
79 => ("00", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "00", "01", "00", "11", "01", "00", "00", "01", "11", "11", "00", "01", "01", "11", "00", "11", "00", "00", "01", "00", "01"),
80 => ("00", "11", "01", "11", "11", "00", "11", "01", "00", "01", "00", "01", "01", "00", "01", "11", "01", "11", "00", "01", "01", "11", "01", "01", "11", "11", "00", "01", "00", "01", "01", "00"),
81 => ("00", "11", "11", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "01", "01", "00", "11", "01", "00", "01", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11"),
82 => ("01", "11", "11", "01", "01", "11", "00", "11", "11", "01", "11", "00", "11", "01", "01", "00", "00", "01", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "00", "01", "00", "01"),
83 => ("01", "01", "01", "11", "01", "11", "01", "00", "01", "01", "01", "01", "01", "11", "01", "00", "01", "11", "11", "00", "11", "01", "00", "11", "00", "01", "01", "11", "01", "01", "11", "01"),
84 => ("00", "00", "01", "01", "01", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "11", "11", "01", "00", "11", "01", "11", "11", "01", "01", "01", "00", "00", "00", "01", "00", "00"),
85 => ("00", "01", "01", "01", "11", "01", "01", "01", "00", "11", "11", "11", "01", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "01", "11", "11", "11", "00", "01"),
86 => ("00", "01", "11", "00", "11", "01", "11", "00", "01", "01", "01", "11", "00", "00", "11", "11", "00", "01", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00", "00", "11", "00", "00"),
87 => ("01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "11", "11", "00", "11", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "01", "01", "01", "11"),
88 => ("00", "11", "01", "01", "01", "00", "11", "00", "11", "00", "11", "01", "00", "11", "01", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "01", "00", "01", "11"),
89 => ("00", "00", "00", "00", "00", "00", "01", "11", "11", "11", "00", "01", "01", "00", "00", "00", "11", "01", "11", "01", "00", "00", "11", "01", "01", "00", "00", "00", "11", "01", "11", "01"),
90 => ("01", "00", "00", "01", "11", "11", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "01", "01", "00", "01", "00", "00", "01", "11", "11", "11", "00", "00", "11", "00", "11", "00"),
91 => ("00", "01", "01", "01", "00", "11", "01", "01", "00", "01", "11", "00", "01", "00", "11", "01", "01", "00", "01", "11", "00", "00", "01", "00", "00", "11", "00", "00", "00", "00", "11", "00"),
92 => ("01", "01", "00", "01", "11", "11", "11", "01", "00", "00", "01", "00", "00", "00", "01", "01", "00", "11", "01", "11", "00", "00", "01", "00", "11", "01", "01", "00", "11", "01", "01", "11"),
93 => ("00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01", "01", "11", "11", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "11", "11", "11", "11"),
94 => ("00", "01", "11", "01", "11", "00", "00", "01", "01", "11", "11", "01", "11", "01", "01", "11", "01", "00", "00", "01", "11", "11", "00", "00", "00", "01", "01", "01", "00", "01", "00", "01"),
95 => ("00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "11", "00", "01", "11", "00", "01", "01", "00", "01", "11", "00", "00", "11", "00", "01", "01", "01", "01", "11", "11"),
96 => ("01", "11", "11", "01", "01", "01", "00", "11", "01", "00", "11", "01", "00", "00", "11", "00", "01", "00", "01", "01", "11", "11", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01"),
97 => ("01", "11", "01", "01", "01", "00", "01", "01", "01", "11", "00", "00", "00", "01", "01", "01", "01", "11", "11", "01", "01", "11", "11", "00", "01", "11", "11", "01", "01", "01", "00", "01"),
98 => ("01", "00", "00", "01", "11", "11", "01", "00", "11", "01", "11", "01", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "11", "01"),
99 => ("01", "00", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "00", "11", "11", "01", "01", "00", "01", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "00", "11"),
100 => ("01", "00", "11", "11", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "00", "00", "00", "11", "11", "00", "00", "11", "00", "01", "01", "11", "01", "11", "00"),
101 => ("01", "01", "00", "00", "11", "01", "01", "00", "11", "11", "01", "00", "01", "11", "01", "00", "11", "01", "11", "01", "00", "01", "01", "00", "11", "00", "01", "01", "00", "11", "00", "01"),
102 => ("00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "00", "11", "11", "00", "00", "00", "00", "00", "01", "11", "11", "11", "00", "11", "11", "11", "00", "00", "01", "01", "00", "01"),
103 => ("01", "00", "11", "01", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "11", "11", "11", "11", "00", "01", "00", "00", "00", "00", "01", "01", "11", "11", "01", "00", "01"),
104 => ("00", "11", "00", "11", "01", "11", "00", "01", "00", "00", "00", "11", "01", "01", "11", "00", "00", "01", "00", "11", "01", "11", "00", "01", "01", "01", "01", "11", "00", "00", "01", "01"),
105 => ("00", "01", "11", "01", "01", "11", "00", "11", "00", "00", "01", "11", "01", "01", "00", "11", "00", "11", "01", "00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "11", "01", "00"),
106 => ("01", "00", "01", "00", "01", "01", "11", "00", "00", "01", "01", "00", "00", "11", "01", "11", "11", "00", "01", "11", "11", "01", "01", "11", "11", "00", "01", "01", "00", "01", "00", "00"),
107 => ("01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "00", "11", "01", "11", "11", "00", "00", "01", "01", "11", "00", "01", "11", "00", "11", "11", "00", "01", "01", "01", "01"),
108 => ("00", "01", "11", "01", "01", "00", "11", "01", "11", "01", "00", "00", "11", "00", "01", "11", "11", "00", "01", "00", "11", "11", "01", "01", "01", "11", "01", "01", "00", "01", "01", "00"),
109 => ("01", "01", "00", "00", "00", "01", "11", "11", "11", "00", "01", "11", "00", "01", "01", "00", "11", "00", "11", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "01", "11", "01"),
110 => ("01", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "00", "11", "01", "11", "01", "01", "00", "11", "01", "00", "01", "11", "00", "11", "01", "01", "11", "11"),
111 => ("00", "11", "01", "01", "00", "01", "11", "01", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "01", "11", "00", "01", "01", "11", "01", "11", "11", "00", "01", "00", "11", "11"),
112 => ("00", "00", "01", "11", "01", "00", "01", "11", "11", "11", "11", "11", "01", "01", "00", "11", "01", "00", "01", "00", "00", "11", "00", "01", "01", "00", "01", "01", "01", "01", "11", "00"),
113 => ("01", "00", "11", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "01", "11", "01", "01", "11", "01", "00", "00", "00", "00", "11", "11", "11", "00", "00", "00", "00", "11", "01"),
114 => ("01", "00", "11", "11", "00", "11", "00", "00", "00", "01", "01", "01", "11", "01", "01", "00", "00", "11", "11", "01", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "00", "00"),
115 => ("01", "00", "01", "11", "11", "00", "00", "01", "11", "01", "01", "00", "11", "00", "11", "00", "01", "01", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "00"),
116 => ("01", "00", "11", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "11", "11", "01", "01", "01", "00", "11", "11", "01", "01", "11", "00", "00", "01", "11", "00", "01"),
117 => ("00", "00", "01", "11", "11", "00", "11", "01", "00", "11", "00", "00", "00", "11", "00", "01", "01", "00", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01", "01", "11", "00", "00"),
118 => ("01", "01", "11", "01", "00", "00", "11", "00", "00", "01", "01", "01", "01", "11", "00", "11", "00", "01", "11", "11", "11", "01", "00", "00", "01", "01", "00", "00", "01", "00", "00", "01"),
119 => ("01", "01", "01", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "00", "00", "11", "11", "00", "11", "11", "01", "01", "01", "01", "11", "11", "11", "00", "00", "01"),
120 => ("00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "01", "11", "01", "01", "11", "01", "11", "00", "11", "00", "01", "00", "11", "01", "00", "00", "01", "11", "01", "01", "01", "00"),
121 => ("00", "11", "00", "11", "11", "01", "01", "11", "01", "00", "11", "11", "01", "01", "00", "01", "00", "11", "11", "00", "00", "00", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00"),
122 => ("00", "00", "00", "00", "11", "01", "01", "00", "01", "00", "11", "01", "00", "01", "01", "01", "01", "11", "11", "11", "01", "00", "00", "00", "00", "11", "11", "01", "01", "11", "00", "11"),
123 => ("00", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "00", "11", "00", "01", "00", "11", "01", "11", "00", "11", "00", "01", "11", "00", "00", "01", "11", "00", "00", "00"),
124 => ("01", "01", "00", "00", "11", "00", "01", "01", "11", "00", "01", "11", "00", "01", "01", "01", "11", "00", "11", "00", "11", "00", "01", "00", "00", "01", "01", "00", "00", "01", "01", "11"),
125 => ("01", "00", "00", "11", "01", "01", "11", "01", "00", "11", "01", "11", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "11", "11", "01", "11", "11", "01", "00", "00", "01", "00"),
126 => ("01", "11", "01", "01", "11", "00", "01", "01", "01", "00", "11", "00", "11", "11", "01", "00", "11", "00", "11", "00", "01", "01", "01", "01", "01", "11", "00", "01", "01", "00", "00", "01"),
127 => ("00", "00", "11", "00", "00", "11", "00", "00", "01", "01", "01", "01", "11", "01", "01", "11", "01", "00", "01", "01", "11", "01", "00", "00", "01", "00", "11", "00", "11", "01", "11", "01"),
128 => ("01", "00", "01", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00", "11", "01", "11", "00", "01", "01", "00", "11", "00", "11", "11", "00", "11", "01", "11", "00", "01", "11", "00"),
129 => ("01", "00", "01", "00", "00", "01", "11", "00", "00", "11", "01", "11", "00", "01", "01", "01", "00", "11", "01", "11", "11", "01", "01", "00", "00", "00", "11", "11", "01", "00", "01", "01"),
130 => ("01", "01", "00", "01", "00", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00", "00", "11", "00", "01", "01", "00", "11", "11", "00", "11", "01", "00", "00", "01", "01", "01", "00"),
131 => ("01", "11", "01", "00", "11", "00", "01", "00", "01", "00", "01", "01", "11", "00", "01", "00", "11", "00", "00", "01", "11", "01", "00", "11", "11", "01", "00", "00", "01", "00", "01", "01"),
132 => ("01", "11", "01", "01", "01", "11", "01", "11", "01", "01", "00", "01", "01", "11", "00", "11", "00", "01", "00", "01", "01", "11", "01", "01", "00", "01", "01", "00", "11", "01", "11", "01"),
133 => ("01", "11", "01", "01", "01", "11", "00", "11", "11", "00", "00", "01", "11", "01", "11", "00", "01", "00", "01", "01", "01", "00", "11", "00", "01", "00", "01", "01", "11", "01", "01", "01"),
134 => ("01", "11", "11", "00", "01", "00", "01", "01", "00", "11", "01", "11", "11", "11", "01", "00", "01", "01", "00", "01", "11", "00", "11", "00", "00", "00", "00", "00", "01", "01", "00", "11"),
135 => ("00", "11", "00", "11", "00", "00", "11", "00", "11", "01", "11", "01", "00", "11", "00", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "01", "00", "11"),
136 => ("01", "00", "00", "01", "00", "11", "11", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "00", "00", "01", "11", "00", "00", "11", "01", "01", "01", "01", "01", "11", "00", "11"),
137 => ("01", "01", "01", "00", "00", "00", "00", "01", "11", "01", "00", "11", "11", "11", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "01", "01", "11", "00", "00", "11", "01", "00"),
138 => ("00", "01", "01", "11", "01", "01", "11", "00", "11", "01", "11", "11", "01", "01", "01", "01", "01", "11", "00", "11", "00", "11", "01", "01", "00", "01", "00", "11", "01", "01", "01", "01"),
139 => ("00", "01", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "11", "00", "11", "01", "01", "11", "00", "01", "11", "01", "00", "01", "11", "11", "11", "01", "00", "11", "00", "01"),
140 => ("01", "11", "01", "01", "11", "01", "01", "00", "00", "01", "01", "00", "01", "00", "00", "00", "11", "01", "01", "01", "11", "11", "01", "11", "01", "01", "11", "01", "01", "01", "00", "00"),
141 => ("01", "00", "00", "01", "00", "01", "01", "00", "00", "01", "11", "00", "00", "11", "00", "01", "00", "00", "00", "11", "11", "11", "00", "01", "00", "01", "01", "11", "00", "01", "11", "11"),
142 => ("01", "11", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "11", "01", "11", "01", "01", "11", "00", "01", "00", "00", "00", "11", "00", "11", "11", "01", "01"),
143 => ("00", "11", "00", "01", "11", "00", "01", "01", "11", "01", "11", "00", "01", "11", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "11", "00", "01", "01", "11", "00", "11"),
144 => ("00", "01", "00", "00", "00", "01", "00", "11", "11", "01", "11", "11", "11", "01", "00", "00", "11", "00", "11", "00", "01", "01", "00", "00", "01", "11", "00", "00", "01", "01", "01", "11"),
145 => ("00", "00", "01", "11", "00", "01", "00", "00", "01", "11", "01", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "00", "01", "11", "01", "11", "01", "11", "01"),
146 => ("01", "01", "00", "11", "00", "11", "01", "00", "01", "11", "00", "01", "01", "01", "11", "00", "00", "11", "01", "11", "11", "01", "01", "01", "00", "11", "01", "11", "00", "00", "00", "00"),
147 => ("01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "11", "00", "11", "11", "11", "00", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11"),
148 => ("00", "00", "01", "01", "00", "01", "01", "01", "11", "01", "01", "00", "11", "00", "11", "01", "01", "11", "11", "00", "11", "01", "01", "00", "01", "00", "00", "11", "11", "01", "00", "01"),
149 => ("00", "00", "00", "11", "01", "11", "01", "01", "01", "00", "01", "00", "01", "00", "11", "11", "11", "00", "00", "00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "01", "11", "01"),
150 => ("01", "01", "11", "01", "01", "01", "01", "00", "00", "01", "01", "00", "00", "11", "11", "01", "01", "01", "01", "00", "01", "11", "01", "11", "11", "11", "00", "00", "01", "11", "01", "01"),
151 => ("01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "11", "00", "01", "11", "11", "00", "01", "01", "00", "01", "11", "11", "01", "00", "01", "00", "01", "11", "01", "00", "01", "11"),
152 => ("00", "01", "01", "01", "00", "11", "00", "11", "01", "00", "01", "01", "00", "11", "01", "11", "01", "00", "11", "01", "00", "01", "01", "01", "01", "01", "01", "11", "11", "01", "01", "11"),
153 => ("01", "01", "01", "01", "00", "11", "00", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "00", "00", "11", "00", "11", "01", "11", "11", "11", "01", "00", "01", "00", "01", "01"),
154 => ("00", "01", "00", "00", "00", "11", "00", "11", "00", "01", "01", "01", "00", "00", "01", "11", "11", "01", "00", "01", "01", "00", "01", "00", "11", "01", "11", "01", "00", "00", "00", "11"),
155 => ("01", "00", "11", "01", "01", "11", "01", "00", "11", "01", "01", "00", "01", "00", "01", "11", "11", "11", "01", "11", "11", "00", "00", "01", "00", "01", "00", "01", "01", "11", "01", "00"),
156 => ("00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "00", "01", "11", "01", "00", "11", "00", "11", "01", "00", "01", "11", "11", "11", "00", "11"),
157 => ("00", "00", "01", "00", "11", "00", "00", "11", "11", "00", "00", "11", "01", "00", "11", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "01", "11", "11", "01", "01", "01", "00"),
158 => ("01", "01", "01", "11", "00", "01", "00", "11", "11", "00", "00", "01", "01", "01", "11", "00", "01", "11", "00", "00", "00", "00", "11", "01", "11", "00", "00", "11", "00", "01", "11", "00"),
159 => ("00", "01", "00", "01", "01", "00", "01", "11", "00", "00", "11", "11", "00", "01", "11", "00", "11", "11", "01", "01", "01", "11", "01", "00", "11", "01", "11", "00", "00", "01", "00", "00"),
160 => ("01", "00", "01", "11", "11", "11", "01", "00", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "11", "11", "00", "11", "01", "00", "00", "01", "01", "11", "01", "01", "00", "01"),
161 => ("01", "01", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "11", "01", "00", "11", "01", "11", "00", "00", "00", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00", "11"),
162 => ("00", "01", "11", "00", "11", "11", "11", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "01", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "00", "00", "00", "00"),
163 => ("01", "00", "00", "00", "00", "11", "01", "00", "01", "01", "11", "01", "01", "00", "00", "00", "11", "11", "01", "00", "00", "11", "01", "01", "01", "01", "01", "11", "11", "00", "11", "11"),
164 => ("01", "11", "00", "00", "00", "01", "00", "11", "01", "01", "01", "01", "01", "00", "01", "11", "11", "11", "00", "01", "00", "01", "01", "11", "11", "01", "11", "00", "00", "11", "00", "00"),
165 => ("00", "01", "01", "00", "01", "00", "11", "01", "00", "01", "00", "00", "01", "11", "00", "00", "01", "01", "11", "00", "00", "01", "01", "11", "00", "00", "01", "11", "01", "11", "11", "11"),
166 => ("00", "11", "01", "01", "01", "11", "11", "11", "00", "00", "00", "01", "00", "01", "00", "11", "00", "11", "01", "01", "00", "00", "11", "11", "01", "11", "01", "01", "00", "00", "00", "01"),
167 => ("01", "11", "00", "01", "01", "00", "11", "00", "01", "11", "00", "11", "11", "00", "01", "00", "01", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "11", "00", "00", "00", "01"),
168 => ("00", "00", "01", "00", "11", "11", "11", "11", "00", "01", "01", "00", "11", "00", "01", "01", "11", "01", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00"),
169 => ("00", "00", "00", "00", "11", "00", "01", "00", "00", "01", "11", "00", "11", "01", "01", "11", "11", "11", "01", "00", "01", "01", "00", "01", "01", "11", "00", "11", "01", "00", "00", "00"),
170 => ("00", "11", "11", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "00", "11", "01", "00", "00", "00", "01", "00", "01", "11", "01", "11"),
171 => ("00", "00", "01", "01", "11", "01", "11", "01", "11", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "11", "11", "00", "00", "01", "11", "11", "00", "01", "01", "11", "00", "01"),
172 => ("00", "01", "01", "01", "01", "01", "00", "01", "00", "11", "11", "11", "00", "00", "11", "00", "01", "11", "01", "11", "11", "11", "01", "01", "01", "00", "00", "00", "01", "01", "01", "00"),
173 => ("01", "00", "00", "00", "11", "11", "01", "11", "01", "11", "01", "11", "00", "01", "01", "01", "00", "01", "01", "00", "01", "01", "01", "00", "11", "11", "00", "01", "00", "01", "11", "00"),
174 => ("01", "01", "11", "00", "11", "01", "00", "01", "01", "11", "11", "01", "01", "01", "00", "01", "00", "01", "11", "01", "01", "11", "00", "01", "01", "00", "01", "00", "01", "00", "11", "00"),
175 => ("00", "11", "01", "00", "00", "00", "00", "00", "11", "01", "01", "00", "11", "11", "01", "00", "11", "11", "00", "00", "01", "00", "01", "01", "01", "11", "01", "00", "00", "01", "11", "00"),
176 => ("00", "01", "00", "01", "00", "11", "11", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00", "00", "01", "11", "00", "11", "11", "00", "01", "00", "00", "00", "01", "00", "00", "00"),
177 => ("00", "00", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "11", "11", "01", "01", "11", "01", "00", "00", "01", "00", "11", "11", "00", "01", "01", "00", "00", "00", "11", "11"),
178 => ("00", "01", "01", "01", "01", "00", "01", "01", "11", "01", "00", "00", "11", "01", "11", "01", "00", "11", "01", "11", "01", "11", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00"),
179 => ("00", "00", "11", "00", "11", "01", "11", "11", "11", "01", "00", "00", "00", "11", "01", "11", "00", "01", "01", "01", "00", "00", "01", "01", "01", "01", "00", "01", "01", "01", "11", "11"),
180 => ("00", "00", "00", "00", "01", "11", "00", "11", "01", "11", "11", "01", "00", "11", "11", "00", "00", "01", "11", "00", "11", "01", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00"),
181 => ("00", "00", "01", "01", "00", "00", "01", "01", "11", "01", "01", "01", "11", "00", "00", "11", "11", "11", "01", "11", "00", "00", "01", "11", "11", "00", "01", "01", "01", "00", "00", "00"),
182 => ("00", "11", "01", "11", "01", "00", "01", "00", "01", "00", "11", "01", "00", "01", "11", "11", "01", "01", "11", "00", "01", "00", "01", "11", "00", "00", "01", "00", "00", "01", "01", "11"),
183 => ("01", "11", "01", "01", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "11", "00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "11", "01", "01", "11", "01", "01", "11"),
184 => ("01", "11", "01", "01", "11", "00", "01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01", "11", "11", "11", "01", "00", "00", "01", "01", "11", "00", "00"),
185 => ("00", "11", "00", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "00", "11", "01", "00", "01", "11", "11", "01", "00", "00", "00", "01", "00", "11", "01", "11", "11", "11", "01"),
186 => ("01", "00", "00", "01", "11", "00", "01", "11", "00", "00", "00", "11", "01", "00", "01", "01", "00", "11", "11", "11", "01", "00", "00", "01", "00", "00", "01", "11", "11", "01", "01", "00"),
187 => ("00", "01", "01", "00", "11", "00", "01", "11", "00", "00", "11", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "11", "00", "11", "00", "11"),
188 => ("00", "11", "11", "00", "00", "11", "00", "00", "00", "11", "11", "01", "01", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "01", "01", "01", "11", "11", "00", "00", "11", "11"),
189 => ("00", "01", "01", "01", "11", "00", "01", "00", "00", "11", "00", "00", "00", "01", "11", "11", "00", "01", "11", "01", "00", "01", "01", "01", "00", "00", "00", "01", "01", "11", "01", "00"),
190 => ("00", "00", "01", "00", "11", "11", "01", "00", "00", "00", "01", "11", "00", "01", "00", "00", "00", "00", "11", "11", "01", "00", "00", "00", "11", "01", "00", "01", "00", "00", "11", "00"),
191 => ("01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "11", "01", "00", "01", "00", "00", "11", "01", "01", "00", "01", "11", "01", "00", "00", "01", "11", "01", "00", "11", "01", "01"),
192 => ("01", "11", "00", "00", "00", "00", "01", "11", "01", "01", "01", "11", "01", "01", "11", "00", "00", "00", "00", "00", "11", "01", "11", "11", "00", "00", "00", "00", "00", "11", "01", "01"),
193 => ("00", "01", "11", "01", "00", "01", "11", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "01", "00", "00", "00", "01", "11", "00", "11", "11", "00", "00", "01", "00", "00", "11"),
194 => ("01", "11", "11", "11", "00", "01", "00", "01", "01", "00", "00", "01", "01", "11", "00", "01", "11", "01", "01", "01", "00", "01", "11", "01", "00", "11", "00", "01", "00", "11", "01", "00"),
195 => ("00", "11", "01", "00", "00", "01", "11", "00", "01", "11", "11", "00", "00", "00", "11", "00", "01", "01", "01", "00", "00", "01", "00", "11", "01", "11", "00", "11", "01", "11", "00", "00"),
196 => ("00", "11", "01", "00", "00", "01", "11", "00", "11", "01", "11", "01", "00", "01", "01", "00", "11", "01", "01", "01", "11", "11", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00"),
197 => ("01", "00", "11", "00", "00", "00", "01", "01", "00", "00", "01", "01", "00", "11", "01", "11", "00", "01", "00", "11", "11", "11", "01", "11", "00", "00", "00", "01", "11", "00", "01", "01"),
198 => ("00", "01", "01", "00", "01", "00", "01", "01", "00", "11", "01", "11", "01", "01", "01", "00", "00", "00", "00", "11", "11", "11", "11", "00", "01", "11", "01", "01", "11", "00", "00", "01"),
199 => ("00", "11", "01", "00", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "01", "01", "11", "11", "00", "00", "11", "00", "01", "01", "01", "00", "00", "00", "01", "00", "11", "01"),
200 => ("01", "11", "00", "11", "00", "11", "01", "01", "11", "11", "01", "00", "00", "11", "11", "11", "00", "00", "11", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
201 => ("00", "00", "11", "00", "11", "00", "11", "00", "01", "01", "00", "11", "00", "01", "11", "00", "11", "11", "00", "01", "01", "00", "00", "01", "00", "11", "00", "01", "00", "00", "00", "01"),
202 => ("00", "11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "11", "01", "01", "00", "00", "11", "00", "01", "11", "01", "00", "01", "01", "11", "00", "00", "00", "00", "11"),
203 => ("00", "11", "01", "01", "11", "00", "01", "01", "01", "11", "00", "11", "01", "11", "01", "00", "00", "01", "01", "00", "01", "11", "00", "01", "00", "00", "11", "11", "01", "11", "00", "01"),
204 => ("01", "01", "00", "00", "00", "01", "01", "00", "11", "00", "00", "01", "11", "00", "01", "01", "01", "00", "01", "11", "01", "00", "11", "11", "11", "00", "00", "01", "11", "01", "11", "01"),
205 => ("00", "11", "11", "01", "01", "11", "00", "00", "00", "11", "11", "01", "11", "00", "01", "00", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "01", "11", "11", "01", "01", "01"),
206 => ("01", "01", "11", "11", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "11", "11", "00", "01", "11", "11", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01"),
207 => ("00", "00", "00", "01", "01", "00", "11", "11", "00", "01", "11", "01", "00", "11", "00", "11", "00", "00", "00", "00", "00", "11", "00", "11", "01", "11", "01", "00", "00", "11", "00", "00"),
208 => ("01", "01", "11", "00", "11", "01", "00", "11", "11", "11", "00", "00", "01", "01", "01", "01", "00", "00", "01", "00", "11", "00", "01", "01", "01", "11", "00", "00", "00", "01", "11", "11"),
209 => ("01", "01", "00", "01", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "01", "11", "11", "11", "11", "01", "01", "01", "11", "01", "11"),
210 => ("01", "01", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "00", "00", "01", "11", "01", "11", "01", "01", "11", "11", "00", "00", "00", "01", "00", "01", "11", "11"),
211 => ("00", "11", "01", "00", "01", "01", "01", "01", "01", "11", "01", "11", "01", "00", "00", "00", "11", "00", "11", "11", "01", "00", "00", "00", "00", "11", "11", "01", "01", "01", "01", "11"),
212 => ("01", "01", "00", "01", "00", "11", "01", "01", "11", "01", "11", "01", "01", "11", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "11", "00", "01", "01", "00", "00", "11"),
213 => ("01", "00", "11", "11", "11", "00", "01", "01", "01", "11", "11", "01", "01", "11", "00", "01", "01", "01", "01", "00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "00", "01", "00"),
214 => ("01", "00", "01", "01", "00", "01", "01", "00", "11", "00", "00", "11", "01", "00", "01", "00", "01", "00", "00", "00", "11", "01", "00", "11", "00", "11", "01", "01", "11", "00", "00", "01"),
215 => ("01", "00", "01", "11", "11", "01", "11", "11", "11", "01", "00", "11", "00", "00", "01", "01", "11", "01", "01", "01", "00", "00", "01", "00", "00", "00", "00", "11", "00", "01", "00", "00"),
216 => ("00", "11", "00", "11", "11", "00", "00", "00", "01", "01", "01", "01", "11", "00", "00", "00", "00", "01", "00", "01", "11", "00", "11", "00", "00", "00", "00", "00", "11", "01", "00", "00"),
217 => ("00", "00", "01", "01", "00", "01", "00", "11", "00", "00", "11", "01", "01", "00", "01", "01", "11", "00", "00", "00", "00", "00", "11", "01", "01", "01", "01", "11", "00", "11", "01", "01"),
218 => ("00", "11", "01", "01", "00", "00", "11", "00", "11", "01", "11", "00", "01", "01", "00", "01", "01", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "01", "11", "11", "01", "00"),
219 => ("00", "00", "00", "00", "00", "01", "11", "11", "11", "00", "01", "01", "00", "11", "01", "11", "00", "01", "01", "01", "11", "01", "00", "01", "01", "00", "01", "00", "11", "00", "11", "01"),
220 => ("01", "01", "11", "11", "01", "11", "00", "00", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "00", "11", "11", "01", "01", "01", "01", "01", "01", "11", "01", "11", "01", "01"),
221 => ("01", "01", "11", "01", "11", "01", "01", "01", "11", "00", "00", "01", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "11", "11", "00", "11", "00", "00", "00", "01", "00", "01"),
222 => ("00", "11", "01", "11", "00", "00", "01", "01", "11", "11", "01", "11", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "01", "00", "11", "00"),
223 => ("01", "01", "01", "01", "01", "11", "01", "00", "11", "01", "01", "01", "11", "01", "00", "11", "11", "11", "00", "01", "00", "11", "00", "00", "01", "11", "00", "01", "01", "00", "01", "11"),
224 => ("01", "01", "01", "00", "11", "01", "11", "11", "00", "00", "01", "11", "01", "11", "01", "00", "11", "00", "01", "00", "00", "01", "11", "00", "00", "11", "00", "01", "00", "01", "00", "01"),
225 => ("00", "11", "00", "00", "01", "11", "01", "00", "00", "00", "11", "01", "00", "00", "11", "01", "01", "11", "01", "01", "11", "11", "11", "00", "00", "00", "11", "00", "01", "00", "00", "01"),
226 => ("00", "01", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "11", "01", "00", "11", "11", "00", "00", "01", "01", "00", "11", "11", "11", "00", "01", "00", "00", "00", "01"),
227 => ("01", "01", "00", "11", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "11", "11", "00", "11", "01", "01", "01", "11", "01", "00", "01", "00", "00", "11", "11", "01", "01"),
228 => ("01", "01", "01", "01", "01", "00", "11", "00", "01", "01", "11", "01", "01", "00", "00", "11", "00", "11", "00", "11", "00", "11", "11", "00", "01", "00", "00", "11", "01", "01", "11", "01"),
229 => ("01", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "11", "01", "00", "01", "11", "01", "00", "11", "01", "00", "00", "00", "11", "11", "01", "01", "01", "01", "00", "01", "00"),
230 => ("01", "01", "00", "11", "01", "00", "00", "00", "11", "00", "01", "01", "11", "00", "11", "01", "11", "01", "01", "01", "01", "01", "01", "00", "11", "00", "11", "11", "01", "01", "01", "01"),
231 => ("01", "00", "01", "01", "00", "00", "11", "00", "01", "01", "11", "01", "00", "00", "01", "11", "11", "00", "01", "11", "00", "00", "01", "11", "11", "11", "11", "01", "01", "00", "00", "00"),
232 => ("01", "01", "01", "00", "11", "11", "01", "00", "11", "01", "00", "00", "00", "00", "11", "11", "01", "11", "11", "01", "00", "01", "00", "00", "11", "01", "01", "11", "01", "00", "00", "00"),
233 => ("00", "00", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "11", "00", "11", "01", "00", "00", "11", "01", "11", "01", "00", "00", "00", "01", "01", "01"),
234 => ("00", "00", "01", "00", "11", "11", "00", "00", "01", "11", "00", "11", "00", "01", "00", "11", "00", "00", "11", "00", "11", "00", "01", "00", "00", "01", "11", "01", "01", "01", "11", "01"),
235 => ("01", "00", "11", "01", "01", "01", "00", "11", "00", "00", "00", "00", "00", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "11", "01", "11", "00", "01", "01", "11", "11", "01"),
236 => ("01", "00", "01", "00", "11", "00", "11", "00", "11", "00", "01", "11", "11", "01", "11", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "00", "11", "00", "00"),
237 => ("00", "01", "01", "11", "01", "01", "11", "11", "01", "01", "01", "11", "00", "11", "00", "01", "01", "00", "11", "01", "00", "11", "00", "11", "00", "00", "00", "00", "01", "00", "00", "11"),
238 => ("01", "11", "01", "01", "00", "00", "11", "00", "11", "01", "00", "11", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "11", "01", "00", "00", "11"),
239 => ("01", "00", "00", "11", "01", "11", "00", "00", "11", "11", "01", "01", "11", "00", "00", "11", "11", "01", "00", "00", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "01"),
240 => ("01", "01", "01", "01", "01", "11", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "11", "01", "00", "01", "01", "01", "11", "00", "01", "11", "11", "01", "11", "00"),
241 => ("01", "01", "01", "11", "01", "11", "00", "01", "00", "00", "11", "11", "01", "00", "11", "00", "00", "01", "00", "11", "01", "01", "00", "00", "00", "01", "00", "11", "00", "11", "00", "11"),
242 => ("00", "00", "01", "01", "00", "01", "01", "01", "11", "00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "11", "00", "11", "11", "00", "01", "01", "00", "11", "01", "01", "11", "11"),
243 => ("01", "01", "00", "11", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "01", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00"),
244 => ("01", "01", "11", "00", "00", "00", "11", "11", "00", "00", "00", "11", "01", "11", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "00", "01", "00", "00", "00", "11", "00", "11"),
245 => ("00", "11", "11", "01", "01", "01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "11", "00", "00", "01", "11", "11", "00", "01", "00", "00", "11", "01", "00", "11", "01", "01", "01"),
246 => ("01", "01", "00", "00", "01", "00", "00", "11", "01", "01", "11", "00", "00", "01", "01", "00", "11", "01", "01", "11", "11", "11", "01", "11", "00", "01", "00", "01", "01", "11", "00", "00"),
247 => ("00", "11", "11", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "00", "00", "11", "11", "01", "01", "11", "00", "01", "00", "11", "11", "01", "00", "01", "01", "01", "00", "01"),
248 => ("01", "01", "11", "11", "11", "01", "00", "00", "00", "01", "11", "11", "01", "00", "00", "01", "01", "00", "01", "01", "01", "11", "11", "00", "11", "11", "01", "00", "01", "00", "01", "00"),
249 => ("01", "00", "00", "11", "11", "00", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "01", "01", "01", "11", "01", "11", "01", "11", "11", "01", "00", "00", "11", "01", "01", "11"),
250 => ("00", "01", "11", "01", "01", "01", "11", "11", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "01", "11", "01", "00", "00", "01", "00", "01", "11", "11", "01", "00"),
251 => ("00", "00", "00", "01", "01", "11", "01", "00", "00", "11", "11", "00", "01", "01", "01", "01", "11", "01", "01", "11", "01", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "11"),
252 => ("01", "01", "11", "01", "11", "11", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "01", "00", "00", "00", "01", "01", "01", "01", "00", "11", "11", "11", "11", "00", "11", "00"),
253 => ("00", "11", "00", "01", "11", "00", "11", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "11", "11", "00", "00", "11", "00", "00"),
254 => ("00", "00", "00", "11", "01", "01", "00", "01", "01", "00", "00", "00", "00", "11", "11", "11", "00", "00", "11", "11", "00", "00", "00", "11", "01", "11", "00", "01", "01", "01", "01", "00"),
255 => ("01", "01", "00", "01", "11", "11", "00", "11", "00", "01", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "11", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "00"),
256 => ("01", "00", "00", "00", "01", "11", "01", "00", "01", "00", "00", "01", "00", "01", "11", "01", "00", "00", "11", "00", "01", "01", "11", "11", "11", "11", "11", "00", "11", "01", "01", "00"),
257 => ("00", "00", "01", "11", "11", "01", "00", "00", "01", "00", "01", "00", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "11", "01", "00", "11", "00", "11", "00", "00", "00", "11"),
258 => ("01", "01", "11", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "00", "01", "11", "00", "01", "11", "00", "01", "11", "01", "01", "00", "01", "11", "11", "01", "00", "11"),
259 => ("01", "01", "01", "00", "01", "01", "00", "11", "00", "11", "11", "01", "00", "01", "11", "01", "00", "01", "01", "00", "01", "00", "00", "01", "00", "11", "11", "01", "11", "00", "11", "01"),
260 => ("00", "00", "01", "00", "11", "01", "00", "01", "11", "11", "00", "00", "01", "11", "01", "00", "01", "11", "01", "00", "00", "00", "01", "01", "11", "00", "01", "01", "01", "11", "01", "01"),
261 => ("00", "00", "00", "11", "01", "01", "11", "11", "01", "01", "11", "01", "11", "00", "01", "00", "11", "00", "00", "11", "01", "11", "01", "00", "00", "00", "00", "00", "00", "01", "11", "00"),
262 => ("01", "01", "11", "01", "00", "11", "11", "11", "01", "00", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "11", "00", "01", "00", "11", "11", "00", "00", "11", "00", "01", "00"),
263 => ("00", "11", "00", "00", "01", "11", "00", "01", "11", "00", "11", "11", "11", "01", "11", "01", "00", "11", "01", "00", "01", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "01"),
264 => ("00", "01", "00", "11", "11", "00", "11", "11", "01", "01", "00", "00", "00", "00", "11", "11", "00", "00", "01", "11", "01", "01", "01", "00", "00", "01", "01", "01", "00", "00", "01", "11"),
265 => ("00", "11", "00", "11", "00", "11", "01", "01", "01", "01", "11", "01", "01", "11", "00", "00", "00", "01", "00", "00", "11", "00", "11", "00", "01", "01", "00", "00", "00", "11", "01", "01"),
266 => ("01", "01", "00", "01", "00", "00", "00", "11", "01", "00", "00", "11", "00", "11", "01", "00", "11", "00", "00", "11", "01", "11", "00", "01", "01", "01", "01", "00", "11", "00", "11", "00"),
267 => ("00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "00", "11", "00", "00", "11", "11", "00", "00", "01", "01", "11", "01", "01", "00", "00", "11", "00", "01", "01"),
268 => ("00", "01", "01", "00", "11", "01", "11", "00", "00", "00", "11", "01", "01", "11", "11", "11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "01", "11", "00", "00", "00", "11", "00"),
269 => ("00", "01", "01", "01", "01", "11", "11", "00", "11", "01", "00", "11", "01", "11", "00", "11", "01", "00", "00", "11", "01", "00", "01", "00", "01", "11", "01", "01", "00", "00", "00", "11"),
270 => ("01", "11", "11", "11", "01", "01", "00", "01", "00", "00", "01", "00", "11", "01", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "01", "00", "11", "00", "00", "11", "01", "01"),
271 => ("00", "01", "11", "00", "01", "00", "01", "00", "01", "01", "00", "01", "00", "11", "01", "01", "00", "01", "11", "01", "01", "11", "11", "11", "00", "11", "11", "00", "00", "00", "01", "01"),
272 => ("01", "11", "00", "00", "11", "01", "00", "00", "00", "11", "01", "00", "11", "01", "01", "11", "01", "11", "01", "00", "00", "00", "01", "00", "00", "11", "11", "00", "01", "00", "01", "00"),
273 => ("00", "01", "01", "11", "00", "00", "11", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01", "00", "00", "11", "00", "11", "00", "00", "00", "01", "11", "01", "00", "11", "01", "11"),
274 => ("00", "11", "00", "01", "00", "00", "00", "00", "11", "01", "00", "01", "00", "01", "01", "00", "11", "00", "11", "00", "11", "01", "11", "00", "00", "11", "01", "01", "01", "00", "01", "01"),
275 => ("01", "11", "01", "00", "00", "00", "11", "01", "01", "00", "01", "00", "11", "01", "00", "00", "11", "00", "00", "00", "01", "11", "01", "11", "00", "00", "00", "00", "00", "00", "11", "11"),
276 => ("00", "01", "11", "01", "00", "00", "00", "01", "00", "00", "11", "00", "11", "01", "01", "11", "11", "00", "00", "01", "11", "01", "00", "01", "11", "11", "00", "00", "00", "00", "01", "01"),
277 => ("00", "00", "11", "00", "11", "11", "00", "01", "01", "01", "11", "01", "00", "00", "11", "00", "01", "11", "11", "00", "00", "00", "00", "00", "01", "00", "01", "01", "11", "01", "01", "01"),
278 => ("01", "11", "01", "00", "01", "01", "11", "01", "00", "11", "00", "11", "00", "11", "01", "11", "01", "00", "00", "01", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "11"),
279 => ("00", "11", "00", "00", "00", "11", "11", "11", "00", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "01", "11", "01", "00", "00", "00", "11", "01", "11", "01", "01", "11", "00"),
280 => ("01", "11", "01", "11", "11", "00", "11", "00", "11", "11", "01", "01", "01", "00", "01", "01", "01", "01", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "00", "00", "11", "01"),
281 => ("01", "01", "01", "00", "11", "00", "01", "01", "01", "00", "00", "11", "11", "01", "01", "00", "01", "00", "00", "11", "00", "11", "11", "01", "01", "00", "01", "01", "11", "00", "01", "00"),
282 => ("01", "01", "01", "00", "01", "00", "11", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "11", "11", "01", "01", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "01"),
283 => ("00", "11", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "11", "00", "01", "00", "11", "11", "11", "01", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "11", "00"),
284 => ("01", "11", "01", "01", "00", "11", "11", "11", "00", "01", "01", "01", "11", "00", "00", "11", "01", "11", "01", "00", "00", "00", "01", "00", "01", "00", "00", "01", "11", "00", "11", "00"),
285 => ("01", "00", "01", "11", "01", "01", "00", "01", "01", "11", "00", "00", "11", "11", "00", "01", "11", "01", "00", "00", "01", "00", "01", "11", "01", "11", "00", "00", "00", "01", "11", "01"),
286 => ("00", "00", "00", "01", "01", "01", "11", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "01", "11", "11", "01", "11", "11", "01", "11", "11", "01", "00", "00", "01", "00", "11"),
287 => ("01", "11", "01", "00", "01", "01", "11", "01", "01", "00", "01", "11", "11", "00", "00", "00", "11", "01", "01", "00", "01", "01", "01", "11", "00", "00", "11", "11", "01", "00", "00", "11"),
288 => ("01", "11", "01", "11", "00", "00", "01", "01", "00", "01", "00", "01", "11", "01", "00", "00", "00", "11", "00", "11", "11", "00", "01", "00", "01", "11", "11", "11", "00", "00", "00", "00"),
289 => ("00", "11", "00", "01", "00", "00", "01", "00", "00", "11", "01", "00", "00", "11", "01", "11", "00", "00", "01", "11", "00", "11", "00", "01", "11", "11", "01", "11", "00", "01", "01", "01"),
290 => ("01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "01", "00", "01", "11", "11", "01", "11", "00", "11", "01", "01", "00", "00", "00", "00", "01", "01", "00", "00", "11", "11", "01"),
291 => ("01", "00", "11", "01", "11", "11", "11", "01", "01", "01", "01", "01", "00", "11", "01", "01", "11", "00", "00", "00", "00", "11", "01", "11", "00", "01", "01", "00", "00", "00", "01", "01"),
292 => ("01", "01", "01", "11", "00", "00", "00", "11", "01", "00", "01", "01", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "11", "00", "01", "11", "11", "11", "00", "01", "01", "11"),
293 => ("01", "11", "00", "01", "11", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "01", "01", "11", "01", "00", "00", "01", "01", "01", "00", "11", "11", "00", "11", "00"),
294 => ("01", "01", "01", "01", "00", "01", "11", "00", "01", "11", "01", "11", "11", "00", "01", "00", "11", "11", "11", "01", "01", "11", "00", "00", "00", "01", "01", "00", "01", "00", "01", "00"),
295 => ("01", "01", "00", "00", "01", "00", "11", "11", "11", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "11", "11", "11", "01", "00", "01", "00", "00", "11", "00", "11", "00"),
296 => ("01", "01", "00", "01", "01", "01", "00", "01", "01", "11", "01", "00", "11", "00", "11", "11", "01", "11", "00", "00", "11", "11", "01", "11", "01", "00", "01", "01", "00", "01", "00", "01"),
297 => ("01", "01", "00", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00", "11", "11", "01", "00", "11", "00", "11", "11", "00", "00", "01", "00", "11", "01", "00", "01", "11"),
298 => ("01", "11", "01", "01", "00", "11", "01", "00", "00", "11", "11", "11", "01", "11", "01", "00", "01", "11", "01", "01", "01", "00", "01", "00", "00", "00", "01", "11", "00", "01", "00", "11"),
299 => ("01", "00", "11", "11", "01", "01", "01", "00", "01", "00", "00", "00", "11", "00", "01", "11", "11", "00", "01", "00", "00", "11", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00"),
300 => ("00", "01", "01", "00", "01", "11", "01", "01", "11", "00", "11", "01", "01", "01", "01", "00", "00", "00", "11", "00", "01", "00", "01", "11", "00", "11", "00", "11", "00", "01", "00", "01"),
301 => ("01", "01", "00", "00", "00", "11", "11", "11", "11", "01", "11", "11", "00", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "01", "01", "01", "01", "01", "11", "01", "01", "01"),
302 => ("01", "11", "11", "11", "11", "01", "01", "00", "00", "11", "01", "00", "00", "11", "01", "01", "00", "00", "00", "00", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "01", "01"),
303 => ("00", "01", "01", "00", "00", "00", "00", "00", "01", "11", "01", "11", "01", "11", "01", "01", "01", "01", "11", "11", "01", "00", "01", "00", "00", "00", "00", "00", "11", "01", "01", "01"),
304 => ("00", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "01", "00", "01", "01", "00", "00", "11", "00", "01", "11", "11", "01", "11", "11", "11", "01", "11", "00", "00", "01", "00"),
305 => ("00", "01", "11", "00", "01", "00", "01", "00", "11", "01", "01", "11", "00", "00", "11", "01", "11", "01", "11", "00", "00", "00", "11", "01", "00", "01", "00", "00", "11", "01", "00", "01"),
306 => ("01", "11", "00", "00", "01", "01", "01", "11", "01", "01", "00", "11", "01", "00", "00", "00", "00", "00", "11", "00", "01", "11", "01", "11", "11", "00", "00", "11", "11", "00", "01", "00"),
307 => ("00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "00", "00", "11", "11", "01", "01", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "11", "11", "00"),
308 => ("00", "01", "00", "01", "11", "00", "01", "01", "01", "01", "01", "00", "11", "11", "01", "01", "00", "11", "00", "11", "00", "00", "01", "00", "00", "11", "00", "00", "11", "01", "00", "01"),
309 => ("00", "00", "11", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "11", "01", "11", "00", "01", "00", "00", "01", "11", "11", "00", "01", "01"),
310 => ("01", "01", "01", "00", "01", "11", "11", "00", "11", "00", "00", "01", "00", "00", "01", "11", "11", "11", "00", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "00", "11", "00"),
311 => ("00", "11", "00", "01", "01", "00", "11", "11", "00", "00", "00", "00", "00", "00", "11", "01", "00", "00", "01", "11", "01", "11", "00", "00", "11", "00", "00", "01", "01", "00", "01", "00"),
312 => ("00", "00", "00", "11", "11", "11", "00", "00", "00", "00", "11", "00", "00", "00", "00", "01", "00", "01", "00", "01", "11", "00", "00", "00", "00", "11", "11", "00", "01", "11", "00", "00"),
313 => ("00", "11", "00", "00", "11", "00", "11", "00", "01", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "11", "11", "00", "11", "11", "01", "01", "00", "01", "00", "11"),
314 => ("00", "11", "01", "11", "00", "11", "01", "00", "11", "01", "11", "00", "01", "01", "00", "11", "11", "01", "01", "00", "01", "00", "00", "00", "01", "11", "01", "01", "00", "00", "01", "00"),
315 => ("00", "11", "00", "00", "11", "01", "00", "11", "00", "01", "00", "11", "01", "01", "11", "01", "11", "00", "01", "01", "00", "00", "01", "00", "00", "01", "01", "00", "11", "11", "11", "00"),
316 => ("01", "01", "11", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "00", "01", "11", "00", "00", "00", "11", "11", "00", "11", "11", "00", "01", "01", "00", "00", "01", "11"),
317 => ("01", "01", "00", "11", "00", "11", "11", "00", "01", "00", "00", "01", "00", "11", "00", "00", "00", "00", "00", "01", "00", "11", "11", "00", "11", "01", "01", "01", "01", "01", "01", "00"),
318 => ("01", "01", "01", "01", "01", "01", "11", "01", "00", "00", "01", "00", "11", "11", "11", "11", "11", "00", "01", "00", "00", "00", "11", "11", "01", "00", "00", "01", "01", "11", "00", "00"),
319 => ("01", "11", "00", "01", "00", "00", "11", "01", "00", "00", "00", "11", "01", "11", "00", "11", "00", "00", "00", "01", "01", "01", "11", "00", "11", "00", "11", "01", "00", "00", "01", "01"),
320 => ("01", "01", "11", "11", "00", "00", "01", "01", "11", "11", "00", "00", "01", "00", "01", "00", "01", "11", "00", "01", "01", "11", "11", "00", "00", "00", "01", "01", "00", "01", "11", "01"),
321 => ("00", "00", "00", "01", "11", "00", "11", "11", "01", "01", "01", "11", "11", "01", "11", "01", "01", "00", "00", "01", "11", "00", "01", "11", "01", "00", "00", "00", "01", "01", "00", "00"),
322 => ("01", "00", "01", "00", "11", "01", "00", "00", "01", "01", "01", "01", "00", "11", "00", "11", "11", "01", "00", "00", "01", "01", "01", "01", "00", "01", "11", "01", "00", "01", "11", "11"),
323 => ("00", "01", "01", "01", "01", "00", "11", "01", "01", "01", "00", "11", "01", "11", "01", "01", "00", "01", "11", "11", "00", "11", "00", "01", "11", "11", "00", "00", "01", "00", "00", "11"),
324 => ("01", "00", "00", "00", "11", "11", "00", "00", "11", "00", "00", "00", "01", "11", "01", "11", "01", "11", "01", "00", "01", "00", "01", "01", "01", "01", "01", "00", "01", "00", "01", "11"),
325 => ("00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "00", "00", "01", "01", "00", "00", "01", "11", "11", "11", "01", "11", "00", "00", "00", "11", "01", "11", "01", "00", "01", "11"),
326 => ("00", "11", "11", "01", "01", "00", "11", "11", "01", "00", "01", "01", "00", "00", "01", "00", "01", "01", "00", "11", "00", "01", "01", "01", "11", "11", "01", "00", "11", "01", "01", "00"),
327 => ("01", "11", "00", "11", "01", "01", "00", "11", "11", "11", "01", "00", "00", "01", "01", "00", "01", "11", "11", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "11"),
328 => ("00", "01", "11", "00", "11", "11", "00", "11", "01", "01", "01", "11", "01", "11", "00", "01", "11", "11", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00"),
329 => ("01", "01", "00", "11", "11", "00", "00", "01", "11", "11", "00", "11", "00", "11", "01", "01", "11", "00", "01", "00", "01", "01", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01"),
330 => ("00", "11", "01", "00", "01", "01", "11", "00", "00", "11", "01", "00", "11", "11", "01", "11", "01", "00", "01", "00", "00", "00", "00", "01", "01", "00", "11", "11", "01", "01", "01", "11"),
331 => ("00", "01", "00", "01", "01", "01", "00", "00", "11", "00", "11", "00", "11", "01", "00", "00", "11", "11", "00", "00", "01", "11", "01", "01", "01", "11", "01", "01", "00", "11", "00", "00"),
332 => ("01", "00", "01", "11", "11", "01", "11", "00", "00", "11", "00", "00", "11", "11", "00", "00", "00", "00", "01", "01", "00", "01", "01", "01", "00", "00", "01", "01", "01", "11", "01", "01"),
333 => ("01", "00", "00", "11", "01", "11", "11", "01", "01", "00", "00", "00", "01", "01", "00", "00", "01", "01", "01", "11", "01", "00", "00", "00", "01", "00", "01", "11", "01", "01", "01", "00"),
334 => ("00", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01", "01", "11", "11", "00", "01", "00", "00", "00", "11", "11", "00", "00", "11", "01", "00", "01", "11", "00", "00"),
335 => ("01", "11", "00", "01", "00", "00", "01", "11", "01", "01", "11", "11", "00", "11", "11", "00", "00", "01", "01", "01", "01", "01", "01", "11", "01", "01", "11", "00", "11", "01", "01", "00"),
336 => ("01", "01", "01", "00", "01", "11", "00", "11", "01", "01", "01", "11", "11", "00", "01", "01", "00", "00", "01", "01", "11", "01", "00", "00", "01", "01", "00", "11", "00", "00", "11", "11"),
337 => ("00", "01", "00", "01", "00", "01", "11", "01", "00", "11", "00", "11", "01", "01", "00", "00", "01", "11", "01", "11", "11", "00", "00", "00", "11", "00", "01", "01", "01", "00", "01", "11"),
338 => ("01", "00", "11", "01", "01", "00", "11", "00", "00", "01", "00", "01", "11", "00", "01", "11", "00", "01", "01", "11", "01", "01", "11", "01", "11", "01", "01", "11", "00", "11", "01", "00"),
339 => ("01", "01", "11", "01", "11", "00", "01", "01", "11", "01", "01", "00", "01", "11", "00", "11", "11", "01", "11", "01", "00", "01", "00", "11", "00", "00", "00", "01", "01", "00", "01", "01"),
340 => ("00", "11", "11", "00", "01", "01", "00", "11", "01", "00", "01", "11", "00", "01", "11", "00", "01", "01", "01", "11", "00", "01", "01", "01", "00", "01", "00", "01", "11", "11", "01", "11"),
341 => ("01", "11", "11", "11", "01", "01", "00", "00", "00", "00", "00", "01", "11", "00", "00", "11", "01", "01", "00", "00", "11", "01", "11", "01", "00", "00", "01", "01", "01", "11", "01", "00"),
342 => ("00", "00", "00", "11", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "01", "00", "01", "01", "01", "11", "01", "01", "00", "00", "00", "11", "11", "01", "11", "11"),
343 => ("01", "01", "00", "01", "01", "01", "00", "11", "11", "01", "01", "01", "01", "00", "01", "01", "11", "00", "01", "11", "01", "00", "11", "01", "01", "01", "01", "00", "11", "11", "01", "11"),
344 => ("01", "01", "00", "01", "11", "11", "01", "00", "01", "01", "00", "01", "11", "01", "11", "11", "00", "11", "11", "00", "00", "00", "01", "01", "00", "00", "11", "01", "01", "11", "00", "00"),
345 => ("00", "11", "00", "00", "01", "01", "00", "11", "00", "11", "11", "01", "00", "01", "00", "00", "01", "01", "01", "00", "11", "11", "01", "01", "01", "00", "00", "11", "11", "00", "01", "01"),
346 => ("00", "00", "00", "00", "11", "01", "00", "01", "00", "00", "11", "11", "11", "11", "01", "01", "00", "11", "11", "00", "00", "00", "00", "01", "11", "00", "11", "00", "00", "00", "01", "01"),
347 => ("00", "01", "01", "00", "01", "01", "01", "01", "01", "11", "01", "01", "01", "00", "00", "01", "11", "00", "00", "00", "11", "00", "01", "11", "01", "01", "11", "00", "11", "11", "01", "00"),
348 => ("01", "01", "00", "00", "11", "01", "11", "01", "00", "01", "01", "01", "11", "00", "01", "01", "01", "01", "11", "11", "00", "00", "01", "01", "11", "00", "01", "01", "11", "01", "00", "01"),
349 => ("00", "11", "01", "11", "11", "01", "11", "01", "00", "01", "11", "01", "01", "00", "00", "00", "01", "00", "11", "01", "00", "11", "00", "01", "01", "00", "01", "00", "01", "00", "00", "00"),
350 => ("01", "01", "00", "01", "01", "01", "00", "00", "11", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00", "00", "11", "11", "00", "11", "11", "01", "11", "00", "11", "00"),
351 => ("01", "01", "11", "00", "11", "01", "11", "00", "01", "11", "01", "01", "11", "00", "01", "00", "01", "00", "11", "01", "11", "00", "00", "11", "01", "01", "01", "00", "00", "00", "00", "11"),
352 => ("01", "00", "01", "11", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "00", "11", "00", "11", "00", "00", "00", "11", "00", "00", "01", "11", "01"),
353 => ("00", "11", "00", "11", "00", "00", "01", "11", "01", "00", "01", "11", "11", "01", "11", "01", "01", "00", "00", "00", "01", "00", "01", "01", "00", "11", "11", "00", "00", "11", "01", "01"),
354 => ("00", "01", "00", "01", "11", "11", "01", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "11", "11", "11", "01", "00", "01", "00", "01", "00", "00", "01", "01", "11"),
355 => ("01", "11", "00", "01", "01", "01", "11", "01", "00", "00", "11", "11", "01", "01", "00", "01", "00", "00", "01", "11", "11", "00", "00", "00", "00", "00", "01", "11", "01", "00", "11", "01"),
356 => ("00", "00", "00", "01", "00", "00", "00", "01", "01", "11", "01", "11", "01", "11", "11", "11", "00", "11", "00", "00", "00", "01", "11", "01", "01", "00", "01", "00", "01", "01", "00", "01"),
357 => ("00", "00", "00", "00", "00", "11", "00", "11", "01", "01", "00", "00", "01", "00", "00", "00", "11", "00", "11", "01", "11", "11", "11", "00", "01", "00", "01", "01", "01", "00", "00", "01"),
358 => ("01", "00", "00", "00", "11", "11", "01", "01", "01", "11", "00", "11", "01", "01", "01", "11", "01", "01", "01", "11", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "00", "00"),
359 => ("00", "00", "01", "01", "00", "11", "11", "11", "00", "01", "00", "00", "11", "01", "00", "01", "11", "01", "00", "00", "00", "00", "01", "11", "01", "00", "00", "00", "11", "00", "11", "11"),
360 => ("01", "11", "00", "01", "01", "00", "11", "01", "11", "01", "11", "01", "00", "01", "01", "11", "00", "01", "01", "00", "00", "01", "00", "11", "01", "11", "11", "00", "00", "01", "01", "00"),
361 => ("01", "00", "11", "00", "00", "01", "01", "01", "00", "01", "00", "11", "01", "01", "00", "00", "01", "00", "00", "01", "01", "01", "00", "11", "00", "11", "01", "11", "11", "11", "01", "00"),
362 => ("00", "11", "00", "00", "01", "11", "00", "11", "01", "01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "01", "01", "00", "11", "01", "11", "11", "01", "11", "00", "11", "01", "01"),
363 => ("00", "01", "00", "01", "01", "00", "01", "11", "11", "00", "00", "01", "00", "00", "11", "00", "01", "00", "01", "01", "11", "01", "11", "01", "11", "11", "00", "00", "11", "11", "01", "00"),
364 => ("01", "11", "00", "00", "00", "01", "01", "11", "01", "00", "00", "01", "11", "11", "00", "11", "00", "01", "11", "00", "01", "11", "00", "01", "00", "00", "00", "00", "01", "00", "01", "11"),
365 => ("00", "01", "00", "11", "00", "01", "11", "01", "01", "01", "01", "00", "11", "11", "00", "01", "01", "01", "11", "00", "11", "01", "01", "01", "01", "01", "00", "11", "01", "00", "01", "01"),
366 => ("01", "00", "00", "01", "00", "01", "11", "11", "00", "11", "11", "00", "00", "11", "01", "01", "00", "00", "01", "01", "00", "00", "11", "00", "00", "11", "11", "01", "01", "00", "00", "11"),
367 => ("01", "01", "01", "01", "11", "01", "01", "00", "11", "00", "01", "11", "00", "01", "00", "01", "11", "01", "01", "00", "11", "01", "01", "01", "01", "01", "11", "00", "11", "11", "00", "11"),
368 => ("00", "01", "01", "00", "01", "01", "11", "01", "11", "11", "11", "01", "11", "00", "11", "00", "00", "01", "00", "01", "11", "00", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01"),
369 => ("00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "01", "11", "00", "00", "00", "00", "01", "00", "00", "01", "01", "00", "11", "01", "11", "11", "11", "01", "01", "00", "00", "11"),
370 => ("01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "01", "11", "11", "11", "01", "11", "01", "00", "00", "01", "01", "00", "01", "11", "11", "01", "11", "01", "00", "11", "01", "00"),
371 => ("01", "00", "01", "01", "00", "11", "00", "00", "00", "11", "00", "00", "00", "11", "00", "01", "00", "01", "01", "11", "01", "11", "11", "00", "01", "01", "00", "01", "00", "11", "11", "01"),
372 => ("01", "01", "01", "01", "00", "11", "00", "01", "00", "11", "00", "00", "11", "00", "00", "00", "01", "11", "11", "00", "01", "11", "00", "00", "00", "11", "01", "01", "01", "00", "11", "00"),
373 => ("01", "00", "00", "01", "11", "01", "01", "11", "00", "00", "00", "00", "01", "11", "01", "00", "01", "01", "01", "11", "11", "00", "00", "00", "11", "11", "01", "00", "11", "01", "00", "00"),
374 => ("00", "01", "01", "00", "00", "01", "00", "00", "11", "11", "00", "01", "00", "00", "01", "01", "11", "00", "00", "00", "11", "01", "11", "11", "00", "11", "01", "01", "11", "01", "01", "00"),
375 => ("00", "01", "11", "00", "00", "01", "11", "00", "01", "00", "01", "00", "11", "00", "11", "00", "00", "01", "00", "00", "11", "11", "01", "01", "00", "11", "11", "00", "00", "01", "00", "01"),
376 => ("00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "11", "00", "01", "11", "00", "01", "11", "00", "00", "00", "01", "11", "11", "11", "00", "00", "00", "00", "11", "01", "01", "01"),
377 => ("01", "00", "00", "01", "01", "01", "01", "01", "11", "00", "00", "11", "01", "01", "11", "00", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "11", "01", "01", "11"),
378 => ("00", "01", "11", "11", "01", "00", "11", "01", "00", "01", "00", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "11", "11", "11", "00", "00", "01", "01", "00"),
379 => ("01", "00", "00", "01", "00", "01", "11", "11", "01", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "00", "11", "00", "01", "11", "11", "01", "00", "01", "01", "01", "01", "01"),
380 => ("01", "11", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "01", "00", "01", "01", "11", "11", "11", "00", "00", "00", "01", "01", "00", "01", "00", "11", "00", "11"),
381 => ("01", "11", "01", "00", "11", "00", "01", "11", "01", "01", "00", "11", "01", "01", "00", "11", "00", "00", "00", "01", "01", "01", "11", "01", "01", "01", "00", "11", "00", "00", "01", "01"),
382 => ("01", "01", "11", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "11", "11", "01", "11", "01", "11", "01", "11", "00", "01", "00", "00", "00", "00", "01", "01"),
383 => ("00", "00", "00", "00", "00", "00", "00", "01", "11", "00", "01", "00", "11", "01", "01", "00", "11", "01", "00", "00", "01", "11", "00", "01", "11", "01", "00", "00", "01", "01", "11", "00"),
384 => ("00", "00", "01", "01", "11", "01", "00", "11", "01", "00", "00", "00", "01", "00", "01", "00", "11", "01", "01", "11", "01", "00", "01", "00", "11", "11", "01", "01", "11", "11", "00", "00"),
385 => ("00", "11", "11", "01", "01", "00", "11", "01", "11", "01", "00", "01", "11", "01", "00", "00", "00", "11", "11", "01", "00", "00", "01", "01", "11", "00", "00", "11", "00", "00", "01", "01"),
386 => ("01", "00", "00", "00", "00", "11", "00", "00", "00", "00", "11", "00", "01", "00", "00", "11", "00", "00", "01", "11", "00", "11", "01", "11", "01", "11", "00", "00", "01", "01", "01", "01"),
387 => ("00", "00", "01", "01", "00", "01", "01", "00", "00", "00", "01", "01", "11", "11", "11", "00", "11", "00", "00", "00", "11", "00", "11", "11", "11", "01", "01", "01", "01", "00", "01", "01"),
388 => ("00", "01", "00", "00", "01", "11", "01", "00", "11", "01", "01", "00", "11", "11", "11", "11", "11", "01", "01", "00", "11", "00", "00", "00", "00", "01", "01", "00", "11", "00", "00", "00"),
389 => ("00", "00", "01", "00", "11", "01", "01", "01", "01", "11", "01", "11", "11", "01", "01", "00", "11", "00", "00", "00", "11", "01", "11", "01", "01", "01", "01", "11", "00", "11", "00", "01"),
390 => ("01", "00", "01", "11", "00", "11", "00", "11", "00", "01", "00", "01", "00", "00", "01", "11", "11", "01", "01", "11", "01", "11", "11", "00", "01", "11", "01", "00", "00", "01", "01", "01"),
391 => ("00", "01", "00", "01", "01", "11", "11", "01", "01", "11", "11", "01", "00", "01", "01", "00", "11", "01", "00", "11", "01", "00", "00", "11", "00", "11", "00", "01", "01", "01", "00", "00"),
392 => ("00", "11", "11", "00", "00", "00", "11", "00", "00", "00", "00", "11", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01"),
393 => ("01", "01", "01", "00", "01", "00", "11", "01", "00", "11", "00", "00", "01", "00", "00", "01", "11", "01", "01", "11", "01", "01", "00", "01", "11", "11", "00", "11", "11", "01", "00", "00"),
394 => ("00", "00", "01", "01", "00", "11", "00", "00", "00", "11", "01", "11", "00", "01", "00", "11", "11", "01", "11", "01", "01", "01", "11", "01", "11", "01", "01", "00", "00", "11", "00", "00"),
395 => ("01", "11", "11", "01", "01", "11", "00", "01", "01", "11", "01", "00", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "11", "11", "11", "01", "01", "11", "00", "00"),
396 => ("01", "00", "11", "11", "11", "00", "00", "00", "01", "01", "00", "01", "01", "00", "01", "00", "11", "00", "00", "01", "01", "00", "11", "11", "01", "00", "01", "11", "00", "11", "00", "00"),
397 => ("00", "01", "11", "00", "00", "01", "00", "01", "00", "00", "01", "11", "11", "00", "00", "01", "00", "00", "00", "00", "11", "11", "01", "11", "11", "01", "11", "01", "00", "01", "01", "00"),
398 => ("01", "01", "00", "00", "00", "00", "00", "01", "11", "11", "11", "00", "01", "11", "11", "11", "01", "01", "11", "01", "01", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "00"),
399 => ("00", "01", "01", "01", "11", "00", "00", "01", "00", "00", "01", "01", "00", "00", "00", "00", "01", "00", "00", "01", "01", "11", "00", "00", "01", "11", "11", "11", "00", "11", "00", "00"),
400 => ("00", "11", "11", "01", "00", "00", "00", "00", "11", "11", "01", "11", "11", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "01", "01", "01", "11"),
401 => ("01", "01", "11", "11", "01", "01", "00", "11", "11", "11", "01", "00", "00", "01", "01", "00", "01", "11", "00", "00", "00", "01", "00", "01", "11", "00", "11", "01", "00", "01", "01", "01"),
402 => ("01", "00", "01", "00", "11", "00", "00", "00", "01", "11", "01", "11", "11", "01", "01", "01", "11", "01", "11", "01", "00", "00", "00", "01", "11", "00", "00", "00", "00", "01", "01", "11"),
403 => ("01", "00", "00", "11", "00", "01", "11", "00", "00", "00", "11", "11", "11", "00", "00", "00", "11", "00", "00", "11", "11", "01", "00", "00", "01", "00", "11", "01", "01", "00", "01", "01"),
404 => ("00", "00", "01", "11", "01", "01", "01", "01", "11", "01", "00", "11", "00", "11", "00", "00", "01", "00", "11", "00", "11", "00", "01", "01", "00", "01", "00", "11", "11", "00", "00", "00"),
405 => ("00", "01", "00", "11", "11", "00", "00", "01", "00", "00", "11", "11", "01", "00", "00", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "01", "11", "00", "01", "00"),
406 => ("01", "00", "11", "11", "00", "11", "01", "00", "00", "00", "01", "00", "11", "01", "01", "00", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "11", "00", "11", "11"),
407 => ("01", "11", "11", "11", "00", "00", "11", "00", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "00", "00", "01", "00", "01", "00", "01", "00", "01", "01", "00", "00", "11"),
408 => ("00", "11", "00", "11", "00", "01", "00", "11", "00", "00", "01", "01", "00", "00", "01", "00", "11", "11", "00", "01", "00", "00", "00", "11", "01", "01", "00", "00", "11", "01", "01", "11"),
409 => ("00", "00", "11", "11", "00", "11", "00", "00", "00", "00", "11", "00", "00", "01", "11", "00", "01", "01", "00", "00", "00", "00", "01", "11", "11", "11", "00", "00", "01", "00", "01", "00"),
410 => ("01", "00", "01", "00", "01", "01", "01", "01", "00", "11", "01", "01", "11", "01", "01", "11", "01", "01", "01", "11", "01", "11", "00", "11", "00", "01", "11", "11", "00", "01", "11", "00"),
411 => ("01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "00", "11", "00", "01", "00", "11", "01", "01", "01", "11", "00", "00", "01", "01", "11", "00", "00", "00", "00", "11", "11", "11"),
412 => ("01", "11", "11", "01", "00", "01", "01", "00", "01", "01", "01", "01", "11", "01", "01", "01", "00", "01", "11", "00", "11", "01", "11", "11", "00", "01", "00", "01", "01", "00", "00", "11"),
413 => ("01", "01", "01", "01", "01", "11", "01", "00", "01", "11", "00", "01", "11", "00", "11", "11", "11", "01", "01", "00", "00", "01", "00", "01", "11", "11", "01", "01", "01", "00", "01", "00"),
414 => ("00", "00", "01", "01", "00", "00", "00", "01", "11", "11", "01", "01", "00", "01", "01", "11", "00", "00", "00", "11", "00", "01", "01", "00", "00", "11", "00", "01", "11", "11", "01", "00"),
415 => ("01", "00", "00", "11", "11", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "11", "01", "00", "01", "00", "00", "11", "01", "01", "01", "01", "00", "11", "00", "11", "11", "11"),
416 => ("00", "01", "00", "00", "11", "11", "11", "01", "11", "11", "11", "00", "01", "00", "00", "01", "01", "01", "11", "01", "11", "01", "11", "01", "01", "01", "00", "01", "01", "00", "01", "00"),
417 => ("01", "11", "00", "11", "01", "01", "01", "01", "00", "01", "11", "01", "01", "01", "00", "11", "01", "00", "11", "01", "00", "00", "00", "11", "00", "01", "00", "01", "01", "00", "01", "11"),
418 => ("01", "01", "00", "01", "11", "01", "00", "11", "01", "11", "00", "00", "01", "01", "11", "00", "00", "01", "11", "11", "11", "01", "11", "00", "00", "01", "01", "01", "00", "01", "01", "01"),
419 => ("01", "11", "00", "01", "11", "00", "01", "01", "11", "01", "01", "00", "01", "00", "11", "11", "11", "01", "00", "11", "01", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "11"),
420 => ("00", "01", "11", "00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "01", "00", "01", "00", "11", "01", "00", "11", "11", "11", "01", "00", "00", "11", "11", "00", "11", "01"),
421 => ("00", "01", "11", "11", "00", "01", "01", "11", "00", "00", "01", "00", "00", "11", "11", "00", "00", "00", "01", "00", "11", "01", "00", "11", "11", "00", "00", "00", "01", "01", "00", "00"),
422 => ("01", "01", "11", "01", "00", "01", "11", "11", "11", "00", "01", "00", "01", "11", "00", "00", "01", "01", "01", "01", "01", "00", "11", "00", "11", "11", "01", "00", "00", "01", "11", "00"),
423 => ("00", "00", "11", "01", "01", "01", "00", "11", "11", "11", "01", "11", "00", "01", "00", "11", "00", "01", "01", "00", "11", "01", "00", "00", "01", "01", "11", "11", "00", "00", "00", "00"),
424 => ("00", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "01", "00", "00", "01", "01", "11", "00", "11", "11", "01", "11", "11", "01", "11", "01"),
425 => ("01", "11", "00", "01", "00", "00", "00", "11", "00", "00", "00", "11", "00", "11", "00", "01", "11", "11", "00", "00", "00", "00", "11", "01", "00", "00", "00", "00", "11", "11", "00", "01"),
426 => ("00", "11", "11", "01", "11", "00", "00", "11", "01", "00", "01", "11", "11", "00", "01", "00", "01", "01", "01", "01", "00", "01", "00", "11", "00", "01", "01", "00", "01", "00", "00", "01"),
427 => ("01", "00", "01", "01", "01", "01", "11", "00", "00", "01", "11", "01", "01", "00", "00", "01", "01", "11", "00", "11", "00", "01", "11", "00", "01", "01", "11", "01", "00", "00", "01", "11"),
428 => ("01", "01", "11", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "00", "01", "00", "01", "01", "01", "11", "01", "01", "01", "11", "01", "00", "01", "11", "00", "11", "11", "01"),
429 => ("00", "00", "00", "00", "01", "00", "11", "01", "11", "00", "11", "01", "01", "01", "01", "01", "01", "11", "00", "01", "00", "00", "01", "00", "01", "00", "00", "01", "00", "01", "01", "00"),
430 => ("00", "00", "00", "01", "11", "01", "01", "00", "01", "01", "01", "11", "01", "11", "11", "01", "00", "01", "01", "11", "11", "00", "11", "00", "00", "01", "01", "01", "00", "00", "01", "01"),
431 => ("01", "11", "11", "00", "01", "00", "11", "11", "01", "11", "01", "01", "01", "01", "11", "00", "01", "01", "01", "00", "00", "00", "00", "11", "00", "01", "00", "11", "11", "00", "00", "00"),
432 => ("01", "00", "01", "01", "11", "11", "00", "01", "00", "01", "01", "11", "01", "01", "11", "01", "00", "01", "00", "01", "11", "11", "01", "00", "00", "11", "00", "01", "11", "00", "00", "01"),
433 => ("00", "00", "00", "01", "11", "01", "00", "01", "01", "00", "00", "00", "00", "11", "11", "11", "01", "00", "01", "01", "11", "00", "01", "11", "01", "00", "00", "11", "01", "00", "01", "01"),
434 => ("01", "01", "00", "01", "11", "11", "11", "01", "01", "11", "01", "00", "00", "00", "01", "01", "11", "01", "01", "00", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "01", "00"),
435 => ("00", "11", "11", "00", "01", "00", "01", "01", "11", "01", "00", "01", "01", "01", "01", "01", "01", "01", "00", "11", "11", "01", "01", "11", "11", "00", "00", "11", "00", "01", "00", "11"),
436 => ("01", "11", "01", "01", "01", "01", "00", "00", "11", "01", "01", "01", "01", "11", "00", "00", "00", "11", "00", "01", "11", "00", "01", "01", "00", "00", "01", "01", "01", "01", "11", "01"),
437 => ("00", "01", "00", "01", "00", "00", "00", "01", "01", "11", "01", "11", "00", "01", "11", "11", "11", "00", "01", "11", "00", "00", "01", "01", "00", "00", "00", "01", "11", "00", "01", "00"),
438 => ("01", "01", "01", "11", "11", "01", "11", "01", "11", "00", "11", "00", "00", "01", "11", "00", "01", "00", "00", "11", "11", "00", "01", "00", "01", "01", "00", "01", "00", "00", "00", "00"),
439 => ("00", "11", "01", "01", "01", "01", "00", "11", "01", "11", "00", "00", "00", "01", "01", "11", "00", "11", "00", "00", "01", "11", "11", "01", "01", "01", "00", "00", "01", "00", "11", "00"),
440 => ("00", "11", "01", "11", "00", "11", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "01", "01", "00", "00", "01", "00", "00", "00", "00", "01", "11", "01", "11", "00", "01", "00"),
441 => ("01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "01", "11", "00", "11", "01", "11", "00", "00", "00", "11", "01", "01", "11", "11", "01", "11", "01", "01", "01", "01", "11", "01"),
442 => ("01", "00", "11", "01", "01", "11", "11", "01", "01", "00", "00", "11", "01", "01", "01", "01", "00", "01", "11", "00", "11", "01", "11", "00", "01", "01", "00", "11", "00", "01", "00", "00"),
443 => ("01", "00", "00", "01", "01", "01", "00", "00", "11", "00", "01", "00", "01", "11", "01", "00", "11", "11", "00", "11", "01", "01", "00", "01", "11", "11", "00", "11", "00", "01", "01", "01"),
444 => ("00", "00", "01", "00", "01", "11", "00", "01", "00", "00", "11", "00", "00", "01", "00", "11", "00", "01", "01", "01", "11", "01", "11", "01", "01", "01", "11", "01", "00", "01", "01", "11"),
445 => ("00", "00", "11", "01", "01", "01", "01", "00", "00", "00", "00", "01", "11", "11", "00", "11", "01", "11", "11", "01", "11", "11", "00", "01", "00", "01", "00", "00", "00", "00", "01", "00"),
446 => ("00", "01", "01", "00", "00", "00", "01", "01", "11", "11", "01", "01", "11", "11", "01", "00", "00", "00", "01", "00", "00", "01", "01", "11", "01", "01", "11", "01", "00", "11", "00", "00"),
447 => ("01", "00", "11", "00", "01", "00", "00", "00", "11", "11", "00", "01", "00", "11", "01", "00", "01", "00", "11", "01", "11", "11", "01", "00", "00", "00", "01", "00", "11", "01", "11", "00"),
448 => ("01", "11", "11", "11", "01", "01", "00", "00", "11", "00", "01", "11", "11", "11", "00", "00", "00", "01", "01", "01", "01", "11", "00", "01", "00", "01", "00", "00", "01", "01", "11", "00"),
449 => ("01", "11", "01", "00", "11", "01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "11", "11", "11", "11", "01", "00", "01", "01", "11", "00", "01", "01", "01", "00", "11", "01", "00"),
450 => ("01", "00", "00", "11", "00", "11", "11", "11", "01", "01", "01", "11", "01", "01", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "01", "11", "01", "00", "00", "01"),
451 => ("01", "11", "00", "11", "01", "11", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "11", "00", "01", "01", "11", "01", "01", "01", "01", "11", "11", "00", "00", "00", "11", "01"),
452 => ("00", "00", "00", "01", "00", "11", "01", "11", "01", "00", "11", "01", "00", "00", "01", "00", "01", "00", "11", "11", "00", "01", "01", "00", "11", "11", "00", "00", "00", "00", "11", "01"),
453 => ("00", "00", "01", "00", "01", "01", "00", "11", "00", "11", "01", "11", "00", "11", "00", "01", "00", "01", "11", "01", "00", "01", "00", "00", "11", "00", "00", "11", "01", "01", "00", "11"),
454 => ("01", "01", "00", "00", "01", "01", "11", "01", "00", "11", "00", "01", "01", "01", "01", "11", "00", "00", "00", "11", "11", "00", "11", "00", "00", "11", "00", "01", "00", "01", "11", "01"),
455 => ("01", "00", "01", "00", "01", "00", "01", "01", "11", "01", "11", "01", "01", "00", "11", "11", "01", "00", "11", "00", "01", "00", "11", "01", "01", "01", "11", "01", "00", "00", "00", "01"),
456 => ("00", "00", "01", "00", "00", "11", "00", "00", "01", "01", "11", "00", "11", "00", "11", "00", "01", "11", "01", "00", "01", "00", "11", "01", "00", "11", "11", "00", "01", "00", "00", "01"),
457 => ("01", "00", "11", "11", "00", "11", "00", "01", "00", "01", "01", "00", "00", "11", "11", "01", "00", "11", "01", "01", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "00", "01"),
458 => ("00", "00", "00", "00", "00", "01", "01", "11", "11", "00", "00", "01", "01", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "01", "01", "00", "11", "01", "11", "00", "00", "11"),
459 => ("00", "11", "01", "01", "01", "11", "01", "11", "00", "01", "01", "00", "01", "00", "01", "11", "00", "01", "00", "01", "11", "11", "00", "00", "01", "01", "00", "00", "01", "11", "11", "01"),
460 => ("01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "00", "11", "11", "11", "01", "11", "00", "01", "11", "00", "00", "00", "01", "00", "11", "01", "00", "00"),
461 => ("00", "00", "00", "01", "00", "01", "00", "11", "01", "00", "01", "00", "11", "01", "11", "00", "01", "00", "11", "11", "00", "00", "00", "01", "11", "00", "01", "01", "01", "01", "11", "11"),
462 => ("01", "11", "11", "01", "01", "00", "01", "00", "11", "00", "00", "00", "11", "00", "11", "00", "01", "01", "01", "01", "11", "11", "11", "00", "00", "00", "00", "01", "01", "01", "11", "01"),
463 => ("00", "01", "01", "01", "11", "11", "00", "11", "00", "00", "00", "01", "00", "00", "01", "01", "01", "11", "01", "11", "01", "00", "11", "00", "01", "11", "00", "01", "11", "00", "01", "00"),
464 => ("00", "01", "11", "00", "00", "00", "00", "00", "00", "11", "01", "11", "01", "01", "00", "11", "00", "00", "11", "01", "00", "00", "01", "11", "01", "01", "00", "00", "00", "00", "00", "01"),
465 => ("00", "00", "00", "11", "01", "01", "01", "01", "01", "11", "01", "01", "01", "01", "00", "00", "00", "01", "01", "01", "01", "11", "00", "11", "11", "00", "00", "01", "11", "01", "11", "00"),
466 => ("00", "11", "01", "00", "01", "11", "00", "00", "01", "11", "00", "11", "00", "00", "01", "11", "00", "01", "00", "01", "00", "00", "11", "00", "00", "01", "01", "00", "00", "00", "11", "00"),
467 => ("00", "01", "01", "01", "01", "01", "01", "01", "11", "01", "01", "11", "11", "01", "00", "11", "00", "01", "11", "11", "01", "00", "11", "01", "01", "00", "00", "01", "00", "11", "00", "11"),
468 => ("00", "00", "00", "11", "01", "00", "00", "00", "01", "01", "01", "11", "11", "01", "11", "11", "01", "11", "00", "00", "01", "01", "01", "01", "00", "11", "00", "01", "00", "01", "00", "11"),
469 => ("00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "00", "01", "00", "11", "01", "11", "01", "01", "00", "11", "00", "00", "00", "00", "00", "11", "01", "00", "11", "11", "11", "00"),
470 => ("01", "01", "11", "11", "11", "00", "00", "00", "11", "01", "00", "00", "01", "11", "00", "11", "00", "00", "01", "01", "01", "11", "01", "01", "01", "01", "01", "00", "00", "01", "00", "00"),
471 => ("01", "11", "11", "01", "00", "00", "11", "00", "00", "00", "11", "01", "01", "00", "11", "01", "01", "11", "01", "01", "00", "01", "01", "11", "01", "00", "11", "01", "00", "11", "01", "00"),
472 => ("00", "11", "01", "11", "00", "11", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "00", "01", "00", "11", "00", "01", "00", "00", "01", "00", "11", "00", "11", "01", "00", "01"),
473 => ("01", "00", "01", "01", "01", "11", "11", "01", "01", "11", "01", "00", "11", "01", "01", "11", "01", "00", "11", "01", "11", "01", "01", "11", "01", "11", "01", "00", "00", "00", "00", "01"),
474 => ("01", "11", "11", "01", "00", "00", "00", "01", "00", "11", "01", "01", "01", "00", "01", "01", "01", "01", "11", "11", "01", "00", "01", "01", "01", "00", "01", "11", "01", "01", "11", "11"),
475 => ("01", "11", "00", "01", "11", "01", "00", "01", "01", "00", "11", "00", "01", "00", "00", "01", "11", "01", "00", "00", "11", "11", "00", "01", "11", "11", "00", "01", "00", "11", "01", "00"),
476 => ("01", "01", "01", "01", "01", "01", "01", "00", "00", "11", "01", "01", "00", "00", "11", "01", "00", "11", "11", "01", "11", "00", "00", "01", "00", "01", "01", "00", "01", "01", "01", "01"),
477 => ("01", "11", "00", "11", "00", "11", "00", "01", "00", "01", "00", "00", "01", "00", "00", "01", "11", "00", "11", "01", "11", "11", "11", "01", "00", "00", "11", "00", "00", "00", "01", "01"),
478 => ("00", "00", "11", "01", "11", "01", "01", "11", "11", "11", "11", "01", "00", "00", "01", "01", "01", "01", "01", "00", "01", "01", "01", "01", "00", "01", "11", "00", "01", "11", "01", "01"),
479 => ("00", "11", "00", "01", "01", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "11", "01", "01", "11", "11", "11", "00", "00", "00", "01", "11", "00", "00", "11", "01", "01", "11"),
480 => ("00", "01", "00", "11", "11", "11", "01", "01", "01", "00", "11", "00", "01", "01", "11", "01", "11", "00", "01", "01", "01", "01", "01", "00", "00", "01", "11", "00", "00", "01", "00", "00"),
481 => ("00", "11", "00", "01", "00", "11", "01", "00", "01", "01", "11", "00", "01", "11", "01", "11", "01", "11", "01", "00", "01", "01", "11", "00", "00", "01", "01", "01", "11", "01", "11", "00"),
482 => ("01", "01", "11", "01", "00", "00", "01", "00", "01", "00", "01", "00", "00", "11", "11", "11", "01", "11", "01", "01", "11", "00", "01", "01", "00", "11", "11", "00", "01", "00", "11", "01"),
483 => ("01", "11", "01", "00", "11", "00", "00", "11", "00", "01", "00", "00", "00", "01", "01", "01", "00", "01", "01", "01", "00", "01", "11", "11", "11", "00", "11", "01", "00", "00", "11", "01"),
484 => ("01", "01", "11", "01", "00", "01", "01", "01", "11", "00", "00", "11", "01", "01", "01", "01", "00", "11", "00", "01", "00", "00", "11", "00", "00", "01", "01", "01", "00", "11", "01", "11"),
485 => ("01", "01", "01", "01", "00", "01", "11", "01", "01", "11", "00", "01", "00", "01", "01", "00", "00", "00", "11", "01", "00", "11", "01", "11", "00", "00", "01", "00", "01", "01", "11", "11"),
486 => ("01", "01", "01", "00", "11", "00", "00", "00", "11", "00", "00", "11", "01", "01", "01", "00", "01", "11", "11", "01", "11", "00", "00", "00", "11", "01", "01", "01", "01", "11", "01", "01"),
487 => ("01", "01", "01", "11", "01", "11", "00", "01", "11", "11", "00", "00", "01", "00", "11", "00", "11", "00", "01", "01", "01", "00", "00", "11", "01", "00", "11", "01", "00", "01", "01", "01"),
488 => ("00", "00", "01", "00", "01", "11", "00", "01", "00", "01", "01", "11", "01", "11", "00", "11", "00", "00", "01", "11", "11", "00", "01", "00", "11", "11", "01", "01", "01", "01", "00", "00"),
489 => ("00", "11", "01", "01", "11", "11", "00", "01", "00", "00", "11", "01", "00", "01", "01", "01", "11", "00", "00", "11", "00", "00", "00", "01", "01", "00", "00", "00", "11", "01", "11", "11"),
490 => ("01", "00", "00", "00", "11", "00", "00", "11", "00", "01", "11", "01", "00", "00", "01", "00", "01", "01", "00", "00", "11", "01", "00", "01", "01", "11", "11", "00", "11", "01", "11", "00"),
491 => ("00", "01", "00", "01", "01", "11", "00", "01", "00", "00", "00", "11", "11", "00", "01", "00", "11", "00", "00", "01", "01", "01", "11", "01", "11", "01", "00", "11", "01", "00", "11", "01"),
492 => ("00", "01", "00", "01", "01", "00", "00", "11", "11", "11", "01", "00", "01", "01", "00", "00", "00", "11", "11", "01", "01", "00", "11", "01", "11", "01", "01", "00", "01", "01", "00", "01"),
493 => ("00", "01", "01", "01", "01", "01", "01", "01", "11", "11", "00", "01", "11", "00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "11", "01", "01", "11", "11", "00", "01"),
494 => ("01", "01", "11", "01", "01", "11", "11", "00", "01", "00", "11", "00", "00", "00", "11", "01", "00", "01", "11", "01", "00", "00", "00", "01", "11", "00", "00", "11", "01", "00", "01", "00"),
495 => ("00", "00", "00", "11", "11", "00", "01", "00", "01", "01", "11", "01", "11", "00", "00", "00", "01", "00", "11", "00", "00", "01", "00", "00", "00", "01", "11", "00", "00", "01", "00", "11"),
496 => ("00", "00", "01", "11", "01", "00", "01", "00", "01", "11", "01", "00", "11", "00", "11", "01", "01", "00", "01", "11", "00", "00", "11", "00", "01", "01", "00", "00", "01", "11", "11", "01"),
497 => ("01", "11", "00", "00", "11", "00", "01", "11", "00", "11", "01", "01", "01", "01", "01", "01", "01", "00", "11", "01", "00", "00", "01", "00", "11", "11", "01", "11", "00", "00", "01", "00"),
498 => ("00", "01", "01", "00", "00", "11", "11", "00", "11", "01", "11", "00", "01", "00", "00", "00", "11", "00", "00", "01", "00", "11", "11", "01", "01", "11", "01", "01", "01", "01", "11", "00"),
499 => ("01", "00", "01", "00", "00", "00", "01", "01", "00", "00", "01", "00", "11", "01", "01", "11", "01", "00", "11", "00", "11", "11", "01", "01", "01", "01", "00", "11", "11", "01", "00", "11")));
end data_to_tcam;
package body data_to_tcam is
end data_to_tcam;